magic
tech sky130A
timestamp 1697831380
<< nwell >>
rect 1745 5485 3105 7030
<< poly >>
rect 1310 7385 1360 7395
rect 1310 7355 1320 7385
rect 1350 7355 1360 7385
rect 1310 7345 1360 7355
rect 1280 6925 1330 6935
rect 1280 6895 1290 6925
rect 1320 6895 1330 6925
rect 1280 6885 1330 6895
rect 1225 4490 1275 4500
rect 1225 4460 1235 4490
rect 1265 4460 1275 4490
rect 1225 4450 1275 4460
rect 1835 4090 1885 4100
rect 1575 4060 1845 4090
rect 1875 4060 1885 4090
rect 1575 2760 1610 4060
rect 1835 4050 1885 4060
rect 490 2725 1610 2760
rect 490 2655 540 2725
rect 680 2655 730 2725
rect 1280 20 1330 30
rect 1160 -10 1290 20
rect 1320 -10 1330 20
rect 1280 -20 1330 -10
rect 1445 0 1495 10
rect 1445 -30 1455 0
rect 1485 -30 1495 0
rect 1445 -40 1495 -30
<< polycont >>
rect 1320 7355 1350 7385
rect 1290 6895 1320 6925
rect 1235 4460 1265 4490
rect 1845 4060 1875 4090
rect 1290 -10 1320 20
rect 1455 -30 1485 0
<< locali >>
rect 1310 7385 1360 7395
rect 1310 7355 1320 7385
rect 1350 7355 1360 7385
rect 1310 7345 1360 7355
rect 1765 6980 1795 7005
rect 1280 6925 1330 6935
rect 1280 6895 1290 6925
rect 1320 6915 1645 6925
rect 1320 6895 1650 6915
rect 1280 6885 1330 6895
rect 1640 6890 1650 6895
rect 1225 4490 1275 4500
rect 1225 4460 1235 4490
rect 1265 4460 1625 4490
rect 1225 4450 1275 4460
rect 1590 4025 1625 4460
rect 1840 4100 1880 4205
rect 1835 4090 1885 4100
rect 1835 4060 1845 4090
rect 1875 4060 1885 4090
rect 1835 4050 1885 4060
rect 1590 3985 1735 4025
rect 1405 2990 1690 3020
rect 1405 90 1435 2990
rect 1665 1525 1670 1570
rect 1155 60 1435 90
rect 1280 20 1330 30
rect 1280 -10 1290 20
rect 1320 -10 1330 20
rect 1280 -20 1330 -10
rect 1445 0 1495 10
rect 1645 0 1675 105
rect 1800 5 1835 10
rect 1445 -30 1455 0
rect 1485 -30 1675 0
rect 1445 -40 1495 -30
<< viali >>
rect 1320 7355 1350 7385
rect 1290 6895 1320 6925
rect 1290 -10 1320 20
rect 1455 -30 1485 0
<< metal1 >>
rect 1310 7385 1495 7395
rect 1310 7355 1320 7385
rect 1350 7355 1495 7385
rect 1310 7345 1495 7355
rect 1280 6925 1330 6935
rect 1280 6895 1290 6925
rect 1320 6895 1330 6925
rect 1280 20 1330 6895
rect 1280 -10 1290 20
rect 1320 -10 1330 20
rect 1280 -20 1330 -10
rect 1445 0 1495 7345
rect 1835 4050 1885 4100
rect 1445 -30 1455 0
rect 1485 -30 1495 0
rect 1445 -40 1495 -30
use bias_generator  bias_generator_0
timestamp 1697827976
transform 1 0 4755 0 1 -45
box -3265 45 -1525 7075
use diffamp  diffamp_0
timestamp 1697750532
transform 1 0 700 0 -1 1340
box -775 -6060 680 1350
<< end >>
