magic
tech sky130A
timestamp 1694482748
<< nwell >>
rect -385 220 -40 360
<< nmos >>
rect -255 80 -240 180
rect -185 80 -170 180
<< pmos >>
rect -255 240 -240 340
rect -185 240 -170 340
<< ndiff >>
rect -310 165 -255 180
rect -310 90 -295 165
rect -270 90 -255 165
rect -310 80 -255 90
rect -240 80 -185 180
rect -170 165 -115 180
rect -170 90 -155 165
rect -130 90 -115 165
rect -170 80 -115 90
<< pdiff >>
rect -310 330 -255 340
rect -310 255 -295 330
rect -270 255 -255 330
rect -310 240 -255 255
rect -240 330 -185 340
rect -240 255 -225 330
rect -200 255 -185 330
rect -240 240 -185 255
rect -170 330 -115 340
rect -170 255 -155 330
rect -130 255 -115 330
rect -170 240 -115 255
<< ndiffc >>
rect -295 90 -270 165
rect -155 90 -130 165
<< pdiffc >>
rect -295 255 -270 330
rect -225 255 -200 330
rect -155 255 -130 330
<< psubdiff >>
rect -365 165 -310 180
rect -365 90 -350 165
rect -325 90 -310 165
rect -365 80 -310 90
<< nsubdiff >>
rect -365 330 -310 340
rect -365 255 -350 330
rect -325 255 -310 330
rect -365 240 -310 255
rect -115 330 -60 340
rect -115 255 -100 330
rect -75 255 -60 330
rect -115 240 -60 255
<< psubdiffcont >>
rect -350 90 -325 165
<< nsubdiffcont >>
rect -350 255 -325 330
rect -100 255 -75 330
<< poly >>
rect -255 340 -240 360
rect -185 340 -170 360
rect -255 180 -240 240
rect -185 180 -170 240
rect -255 60 -240 80
rect -185 60 -170 80
rect -285 50 -240 60
rect -285 25 -275 50
rect -250 25 -240 50
rect -285 15 -240 25
rect -210 50 -165 60
rect -210 25 -200 50
rect -175 25 -165 50
rect -210 15 -165 25
<< polycont >>
rect -275 25 -250 50
rect -200 25 -175 50
<< locali >>
rect -360 330 -260 340
rect -360 255 -350 330
rect -325 255 -295 330
rect -270 255 -260 330
rect -360 245 -260 255
rect -235 330 -190 340
rect -235 255 -225 330
rect -200 255 -190 330
rect -235 245 -190 255
rect -165 330 -65 340
rect -165 255 -155 330
rect -130 255 -100 330
rect -75 255 -65 330
rect -165 245 -65 255
rect -210 215 -190 245
rect -210 195 -145 215
rect -165 175 -145 195
rect -360 165 -260 175
rect -360 90 -350 165
rect -325 90 -295 165
rect -270 90 -260 165
rect -360 80 -260 90
rect -165 165 -120 175
rect -165 90 -155 165
rect -130 90 -120 165
rect -165 80 -120 90
rect -140 60 -120 80
rect -385 50 -240 60
rect -385 40 -275 50
rect -285 25 -275 40
rect -250 25 -240 50
rect -285 15 -240 25
rect -210 50 -165 60
rect -210 25 -200 50
rect -175 25 -165 50
rect -140 40 -40 60
rect -210 15 -165 25
rect -210 -5 -190 15
rect -385 -25 -190 -5
<< viali >>
rect -350 255 -325 330
rect -295 255 -270 330
rect -155 255 -130 330
rect -100 255 -75 330
rect -350 90 -325 165
rect -295 90 -270 165
<< metal1 >>
rect -385 330 -40 340
rect -385 255 -350 330
rect -325 255 -295 330
rect -270 255 -155 330
rect -130 255 -100 330
rect -75 255 -40 330
rect -385 245 -40 255
rect -385 165 -40 175
rect -385 90 -350 165
rect -325 90 -295 165
rect -270 90 -40 165
rect -385 80 -40 90
<< labels >>
rlabel locali -40 50 -40 50 3 Y
port 3 e
rlabel locali -385 -15 -385 -15 7 B
port 1 w
rlabel locali -385 50 -385 50 7 A
port 2 w
rlabel metal1 -385 125 -385 125 7 VN
port 4 w
rlabel metal1 -385 295 -385 295 7 VP
port 5 w
<< end >>
