magic
tech sky130A
timestamp 1697403923
<< nmos >>
rect -510 -40 -460 1160
rect -410 -40 -360 1160
rect -210 -40 -160 1160
rect -20 -40 30 1160
rect 180 -40 230 1160
rect 280 -40 330 1160
rect -510 -1290 -460 -90
rect -410 -1290 -360 -90
rect -210 -1290 -160 -90
rect -20 -1290 30 -90
rect 180 -1290 230 -90
rect 280 -1290 330 -90
rect -610 -2750 -560 -1550
rect -510 -2750 -460 -1550
rect -310 -2750 -260 -1550
rect 80 -2750 130 -1550
rect 280 -2750 330 -1550
rect 380 -2750 430 -1550
rect -715 -3050 485 -3000
rect -715 -3275 485 -3225
rect -385 -4670 -335 -3470
rect -285 -4670 -235 -3470
rect -210 -4670 -160 -3470
rect -20 -4670 30 -3470
rect 55 -4670 105 -3470
rect 155 -4670 205 -3470
rect -385 -5920 -335 -4720
rect -285 -5920 -235 -4720
rect -210 -5920 -160 -4720
rect -20 -5920 30 -4720
rect 55 -5920 105 -4720
rect 155 -5920 205 -4720
<< ndiff >>
rect -560 1150 -510 1160
rect -560 -30 -550 1150
rect -520 -30 -510 1150
rect -560 -40 -510 -30
rect -460 1150 -410 1160
rect -460 -30 -450 1150
rect -420 -30 -410 1150
rect -460 -40 -410 -30
rect -360 1150 -210 1160
rect -360 -30 -350 1150
rect -320 -30 -210 1150
rect -360 -40 -210 -30
rect -160 1150 -20 1160
rect -160 -30 -105 1150
rect -75 -30 -20 1150
rect -160 -40 -20 -30
rect 30 1150 180 1160
rect 30 -30 140 1150
rect 170 -30 180 1150
rect 30 -40 180 -30
rect 230 1150 280 1160
rect 230 -30 240 1150
rect 270 -30 280 1150
rect 230 -40 280 -30
rect 330 1150 380 1160
rect 330 -30 340 1150
rect 370 -30 380 1150
rect 330 -40 380 -30
rect -560 -100 -510 -90
rect -560 -1280 -550 -100
rect -520 -1280 -510 -100
rect -560 -1290 -510 -1280
rect -460 -100 -410 -90
rect -460 -1280 -450 -100
rect -420 -1280 -410 -100
rect -460 -1290 -410 -1280
rect -360 -100 -210 -90
rect -360 -1280 -250 -100
rect -220 -1280 -210 -100
rect -360 -1290 -210 -1280
rect -160 -100 -110 -90
rect -160 -1280 -150 -100
rect -120 -1280 -110 -100
rect -160 -1290 -110 -1280
rect -70 -100 -20 -90
rect -70 -1280 -60 -100
rect -30 -1280 -20 -100
rect -70 -1290 -20 -1280
rect 30 -100 180 -90
rect 30 -1280 40 -100
rect 70 -1280 180 -100
rect 30 -1290 180 -1280
rect 230 -100 280 -90
rect 230 -1280 240 -100
rect 270 -1280 280 -100
rect 230 -1290 280 -1280
rect 330 -100 380 -90
rect 330 -1280 340 -100
rect 370 -1280 380 -100
rect 330 -1290 380 -1280
rect -660 -1560 -610 -1550
rect -660 -2740 -650 -1560
rect -620 -2740 -610 -1560
rect -660 -2750 -610 -2740
rect -560 -1560 -510 -1550
rect -560 -2740 -550 -1560
rect -520 -2740 -510 -1560
rect -560 -2750 -510 -2740
rect -460 -1560 -310 -1550
rect -460 -2740 -450 -1560
rect -420 -2740 -310 -1560
rect -460 -2750 -310 -2740
rect -260 -1560 -210 -1550
rect -260 -2740 -250 -1560
rect -220 -2740 -210 -1560
rect -260 -2750 -210 -2740
rect 30 -1560 80 -1550
rect 30 -2740 40 -1560
rect 70 -2740 80 -1560
rect 30 -2750 80 -2740
rect 130 -1560 280 -1550
rect 130 -2740 240 -1560
rect 270 -2740 280 -1560
rect 130 -2750 280 -2740
rect 330 -1560 380 -1550
rect 330 -2740 340 -1560
rect 370 -2740 380 -1560
rect 330 -2750 380 -2740
rect 430 -1560 480 -1550
rect 430 -2740 440 -1560
rect 470 -2740 480 -1560
rect 430 -2750 480 -2740
rect -715 -2955 485 -2945
rect -715 -2990 25 -2955
rect 475 -2990 485 -2955
rect -715 -3000 485 -2990
rect -715 -3060 485 -3050
rect -715 -3095 25 -3060
rect 475 -3095 485 -3060
rect -715 -3105 485 -3095
rect -715 -3180 485 -3170
rect -715 -3215 -705 -3180
rect -255 -3215 485 -3180
rect -715 -3225 485 -3215
rect -715 -3285 485 -3275
rect -715 -3320 -705 -3285
rect -255 -3320 485 -3285
rect -715 -3330 485 -3320
rect -435 -3480 -385 -3470
rect -435 -4660 -425 -3480
rect -395 -4660 -385 -3480
rect -435 -4670 -385 -4660
rect -335 -3480 -285 -3470
rect -335 -4660 -325 -3480
rect -295 -4660 -285 -3480
rect -335 -4670 -285 -4660
rect -235 -4670 -210 -3470
rect -160 -3480 -110 -3470
rect -160 -4660 -150 -3480
rect -120 -4660 -110 -3480
rect -160 -4670 -110 -4660
rect -70 -3480 -20 -3470
rect -70 -4660 -60 -3480
rect -30 -4660 -20 -3480
rect -70 -4670 -20 -4660
rect 30 -4670 55 -3470
rect 105 -3480 155 -3470
rect 105 -4660 115 -3480
rect 145 -4660 155 -3480
rect 105 -4670 155 -4660
rect 205 -3480 255 -3470
rect 205 -4660 215 -3480
rect 245 -4660 255 -3480
rect 205 -4670 255 -4660
rect -435 -4730 -385 -4720
rect -435 -5910 -425 -4730
rect -395 -5910 -385 -4730
rect -435 -5920 -385 -5910
rect -335 -4730 -285 -4720
rect -335 -5910 -325 -4730
rect -295 -5910 -285 -4730
rect -335 -5920 -285 -5910
rect -235 -5920 -210 -4720
rect -160 -4735 -20 -4720
rect -160 -5905 -145 -4735
rect -35 -5905 -20 -4735
rect -160 -5920 -20 -5905
rect 30 -5920 55 -4720
rect 105 -4730 155 -4720
rect 105 -5910 115 -4730
rect 145 -5910 155 -4730
rect 105 -5920 155 -5910
rect 205 -4730 255 -4720
rect 205 -5910 215 -4730
rect 245 -5910 255 -4730
rect 205 -5920 255 -5910
<< ndiffc >>
rect -550 -30 -520 1150
rect -450 -30 -420 1150
rect -350 -30 -320 1150
rect -105 -30 -75 1150
rect 140 -30 170 1150
rect 240 -30 270 1150
rect 340 -30 370 1150
rect -550 -1280 -520 -100
rect -450 -1280 -420 -100
rect -250 -1280 -220 -100
rect -150 -1280 -120 -100
rect -60 -1280 -30 -100
rect 40 -1280 70 -100
rect 240 -1280 270 -100
rect 340 -1280 370 -100
rect -650 -2740 -620 -1560
rect -550 -2740 -520 -1560
rect -450 -2740 -420 -1560
rect -250 -2740 -220 -1560
rect 40 -2740 70 -1560
rect 240 -2740 270 -1560
rect 340 -2740 370 -1560
rect 440 -2740 470 -1560
rect 25 -2990 475 -2955
rect 25 -3095 475 -3060
rect -705 -3215 -255 -3180
rect -705 -3320 -255 -3285
rect -425 -4660 -395 -3480
rect -325 -4660 -295 -3480
rect -150 -4660 -120 -3480
rect -60 -4660 -30 -3480
rect 115 -4660 145 -3480
rect 215 -4660 245 -3480
rect -425 -5910 -395 -4730
rect -325 -5910 -295 -4730
rect -145 -5905 -35 -4735
rect 115 -5910 145 -4730
rect 215 -5910 245 -4730
<< psubdiff >>
rect -610 1145 -560 1160
rect -610 -25 -595 1145
rect -575 -25 -560 1145
rect -610 -40 -560 -25
rect 380 1145 430 1160
rect 380 -25 395 1145
rect 415 -25 430 1145
rect 380 -40 430 -25
rect -610 -105 -560 -90
rect -610 -1275 -595 -105
rect -575 -1275 -560 -105
rect -610 -1290 -560 -1275
rect 380 -105 430 -90
rect 380 -1275 395 -105
rect 415 -1275 430 -105
rect 380 -1290 430 -1275
rect -485 -3485 -435 -3470
rect -485 -4655 -470 -3485
rect -450 -4655 -435 -3485
rect -485 -4670 -435 -4655
rect 255 -3485 305 -3470
rect 255 -4655 270 -3485
rect 290 -4655 305 -3485
rect 255 -4670 305 -4655
<< psubdiffcont >>
rect -595 -25 -575 1145
rect 395 -25 415 1145
rect -595 -1275 -575 -105
rect 395 -1275 415 -105
rect -470 -4655 -450 -3485
rect 270 -4655 290 -3485
<< poly >>
rect 0 1320 460 1350
rect 0 1230 30 1320
rect -510 1220 -460 1230
rect -510 1190 -500 1220
rect -470 1190 -460 1220
rect -510 1160 -460 1190
rect -410 1220 -360 1230
rect -410 1190 -400 1220
rect -370 1190 -360 1220
rect -410 1160 -360 1190
rect -210 1185 30 1230
rect -210 1160 -160 1185
rect -20 1160 30 1185
rect 180 1220 230 1230
rect 180 1190 190 1220
rect 220 1190 230 1220
rect 180 1160 230 1190
rect 280 1220 330 1230
rect 280 1190 290 1220
rect 320 1190 330 1220
rect 280 1160 330 1190
rect -510 -90 -460 -40
rect -410 -90 -360 -40
rect -210 -90 -160 -40
rect -20 -90 30 -40
rect 180 -90 230 -40
rect 280 -90 330 -40
rect -510 -1320 -460 -1290
rect -410 -1315 -360 -1290
rect -210 -1315 -160 -1290
rect -20 -1315 30 -1290
rect 180 -1315 230 -1290
rect -510 -1350 -500 -1320
rect -470 -1350 -460 -1320
rect -510 -1360 -460 -1350
rect 280 -1320 330 -1290
rect 280 -1350 290 -1320
rect 320 -1350 330 -1320
rect 280 -1360 330 -1350
rect -310 -1495 640 -1445
rect -610 -1550 -560 -1535
rect -510 -1550 -460 -1535
rect -310 -1550 -260 -1495
rect 80 -1550 130 -1495
rect 280 -1550 330 -1535
rect 380 -1550 430 -1535
rect -610 -2780 -560 -2750
rect -610 -2810 -600 -2780
rect -570 -2810 -560 -2780
rect -610 -2820 -560 -2810
rect -510 -2845 -460 -2750
rect -310 -2775 -260 -2750
rect 80 -2775 130 -2750
rect 280 -2845 330 -2750
rect 380 -2780 430 -2750
rect 380 -2810 390 -2780
rect 420 -2810 430 -2780
rect 380 -2820 430 -2810
rect -510 -2895 680 -2845
rect -730 -3050 -715 -3000
rect 485 -3050 570 -3000
rect 515 -3225 570 -3050
rect -730 -3275 -715 -3225
rect 485 -3275 570 -3225
rect -285 -3385 -160 -3375
rect -435 -3415 -335 -3405
rect -435 -3445 -425 -3415
rect -395 -3445 -335 -3415
rect -435 -3455 -335 -3445
rect -385 -3470 -335 -3455
rect -285 -3415 -200 -3385
rect -170 -3415 -160 -3385
rect -285 -3425 -160 -3415
rect -20 -3385 105 -3375
rect -20 -3415 -10 -3385
rect 20 -3415 105 -3385
rect -20 -3425 105 -3415
rect -285 -3470 -235 -3425
rect -210 -3470 -160 -3450
rect -20 -3470 30 -3450
rect 55 -3470 105 -3425
rect 155 -3415 255 -3405
rect 155 -3445 215 -3415
rect 245 -3445 255 -3415
rect 155 -3455 255 -3445
rect 155 -3470 205 -3455
rect -385 -4720 -335 -4670
rect -285 -4720 -235 -4670
rect -210 -4720 -160 -4670
rect -20 -4720 30 -4670
rect 55 -4720 105 -4670
rect 155 -4720 205 -4670
rect -385 -5945 -335 -5920
rect -385 -5975 -375 -5945
rect -345 -5975 -335 -5945
rect -385 -5985 -335 -5975
rect -285 -5945 -235 -5920
rect -210 -5935 -160 -5920
rect -285 -5975 -275 -5945
rect -245 -5975 -235 -5945
rect -285 -5985 -235 -5975
rect -20 -6020 30 -5920
rect 55 -5945 105 -5920
rect 55 -5975 65 -5945
rect 95 -5975 105 -5945
rect 55 -5985 105 -5975
rect 155 -5945 205 -5920
rect 155 -5975 165 -5945
rect 195 -5975 205 -5945
rect 155 -5985 205 -5975
rect -20 -6050 610 -6020
<< polycont >>
rect -500 1190 -470 1220
rect -400 1190 -370 1220
rect 190 1190 220 1220
rect 290 1190 320 1220
rect -500 -1350 -470 -1320
rect 290 -1350 320 -1320
rect -600 -2810 -570 -2780
rect 390 -2810 420 -2780
rect -425 -3445 -395 -3415
rect -200 -3415 -170 -3385
rect -10 -3415 20 -3385
rect 215 -3445 245 -3415
rect -375 -5975 -345 -5945
rect -275 -5975 -245 -5945
rect 65 -5975 95 -5945
rect 165 -5975 195 -5945
<< locali >>
rect 190 1250 460 1280
rect 190 1230 220 1250
rect -510 1220 -460 1230
rect -510 1215 -500 1220
rect -555 1190 -500 1215
rect -470 1190 -460 1220
rect -555 1180 -460 1190
rect -410 1220 -360 1230
rect -410 1190 -400 1220
rect -370 1190 -360 1220
rect -410 1180 -360 1190
rect 180 1220 230 1230
rect 180 1190 190 1220
rect 220 1190 230 1220
rect 180 1180 230 1190
rect 280 1220 330 1230
rect 280 1190 290 1220
rect 320 1215 330 1220
rect 320 1190 375 1215
rect 280 1180 375 1190
rect -555 1160 -515 1180
rect 335 1160 375 1180
rect -610 1150 -510 1160
rect -610 1145 -550 1150
rect -610 -25 -595 1145
rect -575 -25 -550 1145
rect -610 -30 -550 -25
rect -520 -30 -510 1150
rect -610 -40 -510 -30
rect -460 1150 -410 1160
rect -460 -30 -450 1150
rect -420 -30 -410 1150
rect -460 -40 -410 -30
rect -360 1150 -310 1160
rect -360 -30 -350 1150
rect -320 -30 -310 1150
rect -360 -40 -310 -30
rect -115 1150 -65 1155
rect -115 -30 -105 1150
rect -75 -30 -65 1150
rect -115 -40 -65 -30
rect 130 1150 180 1160
rect 130 -30 140 1150
rect 170 -30 180 1150
rect 130 -40 180 -30
rect 230 1150 280 1160
rect 230 -30 240 1150
rect 270 -30 280 1150
rect 230 -40 280 -30
rect 330 1150 430 1160
rect 330 -30 340 1150
rect 370 1145 430 1150
rect 370 -25 395 1145
rect 415 -25 430 1145
rect 370 -30 430 -25
rect 330 -40 430 -30
rect -610 -100 -510 -90
rect -450 -95 -420 -40
rect -610 -105 -550 -100
rect -610 -1275 -595 -105
rect -575 -1275 -550 -105
rect -610 -1280 -550 -1275
rect -520 -1280 -510 -100
rect -610 -1290 -510 -1280
rect -460 -100 -410 -95
rect -460 -1280 -450 -100
rect -420 -1280 -410 -100
rect -460 -1290 -410 -1280
rect -555 -1310 -515 -1290
rect -555 -1320 -460 -1310
rect -555 -1340 -500 -1320
rect -510 -1350 -500 -1340
rect -470 -1350 -460 -1320
rect -510 -1360 -460 -1350
rect -350 -1405 -320 -40
rect -260 -100 -210 -95
rect -260 -1280 -250 -100
rect -220 -1280 -210 -100
rect -260 -1290 -210 -1280
rect -160 -100 -110 -95
rect -160 -1280 -150 -100
rect -120 -1280 -110 -100
rect -160 -1290 -110 -1280
rect -70 -100 -20 -95
rect -70 -1280 -60 -100
rect -30 -1280 -20 -100
rect -70 -1290 -20 -1280
rect 30 -100 80 -95
rect 30 -1280 40 -100
rect 70 -1280 80 -100
rect 30 -1290 80 -1280
rect -550 -1435 -320 -1405
rect -550 -1550 -520 -1435
rect -660 -1560 -610 -1550
rect -660 -2740 -650 -1560
rect -620 -2740 -610 -1560
rect -660 -2750 -610 -2740
rect -560 -1560 -510 -1550
rect -560 -2740 -550 -1560
rect -520 -2740 -510 -1560
rect -560 -2750 -510 -2740
rect -460 -1560 -410 -1550
rect -250 -1555 -220 -1290
rect -460 -2740 -450 -1560
rect -420 -2740 -410 -1560
rect -460 -2750 -410 -2740
rect -260 -1560 -210 -1555
rect -260 -2740 -250 -1560
rect -220 -2740 -210 -1560
rect -260 -2750 -210 -2740
rect -655 -2770 -615 -2750
rect -655 -2780 -560 -2770
rect -655 -2805 -600 -2780
rect -610 -2810 -600 -2805
rect -570 -2810 -560 -2780
rect -610 -2820 -560 -2810
rect -450 -3170 -420 -2750
rect -715 -3180 -245 -3170
rect -715 -3215 -705 -3180
rect -255 -3215 -245 -3180
rect -715 -3225 -245 -3215
rect -715 -3285 -245 -3275
rect -715 -3320 -705 -3285
rect -255 -3320 -245 -3285
rect -715 -3330 -245 -3320
rect -435 -3415 -385 -3405
rect -435 -3445 -425 -3415
rect -395 -3445 -385 -3415
rect -435 -3470 -385 -3445
rect -485 -3480 -385 -3470
rect -325 -3475 -295 -3330
rect -150 -3375 -120 -1290
rect -210 -3385 -120 -3375
rect -210 -3415 -200 -3385
rect -170 -3415 -120 -3385
rect -210 -3425 -120 -3415
rect -150 -3470 -120 -3425
rect -60 -3375 -30 -1290
rect 40 -1550 70 -1290
rect 140 -1405 170 -40
rect 240 -95 270 -40
rect 230 -100 280 -95
rect 230 -1280 240 -100
rect 270 -1280 280 -100
rect 230 -1290 280 -1280
rect 330 -100 430 -90
rect 330 -1280 340 -100
rect 370 -105 430 -100
rect 370 -1275 395 -105
rect 415 -1275 430 -105
rect 370 -1280 430 -1275
rect 330 -1290 430 -1280
rect 330 -1310 375 -1290
rect 280 -1320 375 -1310
rect 280 -1350 290 -1320
rect 320 -1340 375 -1320
rect 320 -1350 330 -1340
rect 280 -1360 330 -1350
rect 140 -1435 370 -1405
rect 340 -1550 370 -1435
rect 30 -1560 80 -1550
rect 30 -2740 40 -1560
rect 70 -2740 80 -1560
rect 30 -2750 80 -2740
rect 230 -1560 280 -1550
rect 230 -2740 240 -1560
rect 270 -2740 280 -1560
rect 230 -2750 280 -2740
rect 330 -1560 380 -1550
rect 330 -2740 340 -1560
rect 370 -2740 380 -1560
rect 330 -2750 380 -2740
rect 430 -1560 480 -1550
rect 430 -2740 440 -1560
rect 470 -2740 480 -1560
rect 430 -2750 480 -2740
rect 240 -2945 270 -2750
rect 435 -2770 475 -2750
rect 380 -2780 475 -2770
rect 380 -2810 390 -2780
rect 420 -2805 475 -2780
rect 420 -2810 430 -2805
rect 380 -2820 430 -2810
rect 15 -2955 485 -2945
rect 15 -2990 25 -2955
rect 475 -2990 485 -2955
rect 15 -3000 485 -2990
rect 15 -3060 485 -3050
rect 15 -3095 25 -3060
rect 475 -3095 485 -3060
rect 15 -3105 485 -3095
rect -60 -3385 30 -3375
rect -60 -3415 -10 -3385
rect 20 -3415 30 -3385
rect -60 -3425 30 -3415
rect -60 -3470 -30 -3425
rect -485 -3485 -425 -3480
rect -485 -4655 -470 -3485
rect -450 -4655 -425 -3485
rect -485 -4660 -425 -4655
rect -395 -4660 -385 -3480
rect -485 -4670 -385 -4660
rect -330 -3480 -290 -3475
rect -330 -4660 -325 -3480
rect -295 -4660 -290 -3480
rect -330 -4665 -290 -4660
rect -160 -3480 -110 -3470
rect -160 -4660 -150 -3480
rect -120 -4660 -110 -3480
rect -425 -4725 -395 -4670
rect -325 -4720 -295 -4665
rect -160 -4670 -110 -4660
rect -70 -3480 -20 -3470
rect 115 -3475 145 -3105
rect 205 -3415 255 -3405
rect 205 -3445 215 -3415
rect 245 -3445 255 -3415
rect 205 -3470 255 -3445
rect -70 -4660 -60 -3480
rect -30 -4660 -20 -3480
rect -70 -4670 -20 -4660
rect 110 -3480 150 -3475
rect 110 -4660 115 -3480
rect 145 -4660 150 -3480
rect 110 -4665 150 -4660
rect 205 -3480 305 -3470
rect 205 -4660 215 -3480
rect 245 -3485 305 -3480
rect 245 -4655 270 -3485
rect 290 -4655 305 -3485
rect 245 -4660 305 -4655
rect 115 -4720 145 -4665
rect 205 -4670 305 -4660
rect -430 -4730 -390 -4725
rect -430 -5910 -425 -4730
rect -395 -5910 -390 -4730
rect -430 -5935 -390 -5910
rect -335 -4730 -285 -4720
rect -335 -5910 -325 -4730
rect -295 -5910 -285 -4730
rect -335 -5915 -285 -5910
rect -155 -4730 -25 -4725
rect -155 -4735 -105 -4730
rect -75 -4735 -25 -4730
rect -155 -5905 -145 -4735
rect -35 -5905 -25 -4735
rect -155 -5915 -25 -5905
rect 105 -4730 155 -4720
rect 215 -4725 245 -4670
rect 105 -5910 115 -4730
rect 145 -5910 155 -4730
rect 105 -5915 155 -5910
rect 210 -4730 250 -4725
rect 210 -5910 215 -4730
rect 245 -5910 250 -4730
rect 210 -5935 250 -5910
rect -430 -5945 -335 -5935
rect -430 -5970 -375 -5945
rect -385 -5975 -375 -5970
rect -345 -5975 -335 -5945
rect -385 -5985 -335 -5975
rect -285 -5945 -235 -5935
rect -285 -5975 -275 -5945
rect -245 -5975 -235 -5945
rect -285 -5985 -235 -5975
rect 55 -5945 105 -5935
rect 55 -5975 65 -5945
rect 95 -5975 105 -5945
rect 55 -5985 105 -5975
rect 155 -5945 250 -5935
rect 155 -5975 165 -5945
rect 195 -5970 250 -5945
rect 195 -5975 205 -5970
rect 155 -5985 205 -5975
<< viali >>
rect -400 1190 -370 1220
rect 190 1190 220 1220
rect -550 -30 -520 1150
rect -105 -30 -75 1150
rect 340 -30 370 1150
rect -550 -1280 -520 -100
rect -650 -2740 -620 -1560
rect 340 -1280 370 -100
rect 440 -2740 470 -1560
rect -425 -4660 -395 -3480
rect 215 -4660 245 -3480
rect -425 -5910 -395 -4730
rect -105 -4735 -75 -4730
rect -105 -5900 -75 -4735
rect 215 -5910 245 -4730
rect -275 -5975 -245 -5945
rect 65 -5975 95 -5945
<< metal1 >>
rect -410 1220 -360 1230
rect 180 1220 230 1230
rect -410 1190 -400 1220
rect -370 1190 190 1220
rect 220 1190 230 1220
rect -410 1180 -360 1190
rect 180 1180 230 1190
rect -560 1150 -510 1160
rect -560 -30 -550 1150
rect -520 -30 -510 1150
rect -560 -100 -510 -30
rect -115 1150 -65 1155
rect -115 -30 -105 1150
rect -75 -30 -65 1150
rect -115 -40 -65 -30
rect 330 1150 380 1165
rect 330 -30 340 1150
rect 370 -30 380 1150
rect -560 -1280 -550 -100
rect -520 -1280 -510 -100
rect -560 -1290 -510 -1280
rect -660 -1560 -610 -1550
rect -660 -2740 -650 -1560
rect -620 -2740 -610 -1560
rect -660 -2750 -610 -2740
rect -435 -3480 -385 -3470
rect -435 -4660 -425 -3480
rect -395 -4660 -385 -3480
rect -435 -4730 -385 -4660
rect -105 -4725 -75 -40
rect 330 -100 380 -30
rect 330 -1280 340 -100
rect 370 -1280 380 -100
rect 330 -1285 380 -1280
rect 430 -1560 480 -1550
rect 430 -2740 440 -1560
rect 470 -2740 480 -1560
rect 430 -2750 480 -2740
rect 205 -3480 255 -3470
rect 205 -4660 215 -3480
rect 245 -4660 255 -3480
rect -435 -5910 -425 -4730
rect -395 -5910 -385 -4730
rect -110 -4730 -70 -4725
rect -110 -5900 -105 -4730
rect -75 -5900 -70 -4730
rect -110 -5910 -70 -5900
rect 205 -4730 255 -4660
rect 205 -5910 215 -4730
rect 245 -5910 255 -4730
rect -435 -5920 -385 -5910
rect 205 -5920 255 -5910
rect -285 -5945 -235 -5935
rect -285 -5975 -275 -5945
rect -245 -5955 -235 -5945
rect 55 -5945 105 -5935
rect 55 -5955 65 -5945
rect -245 -5975 65 -5955
rect 95 -5975 105 -5945
rect -285 -5985 105 -5975
<< labels >>
flabel space 825 1060 1035 1270 0 FreeSans 800 0 0 0 dummy
flabel space 825 -1180 1035 -970 0 FreeSans 800 0 0 0 dummy
<< end >>
