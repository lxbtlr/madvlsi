magic
tech sky130A
timestamp 1697163232
<< error_p >>
rect -2845 1515 -2795 2715
rect -2745 1515 -2695 2715
rect -2645 1515 -2620 2715
rect -2570 1515 -2540 2715
rect -2490 1515 -2465 2715
rect -2415 1515 -2385 2715
rect -2335 1515 -2285 2715
rect -2235 1515 -2210 2715
rect -2160 1515 -2135 2715
rect -2085 1515 -2060 2715
rect -2010 1515 -1985 2715
rect -1935 1515 -1885 2715
rect -1835 1515 -1785 2715
rect -3035 -95 -2985 1105
rect -2935 -95 -2885 1105
rect -2835 -95 -2785 1105
rect -2735 -95 -2685 1105
rect -2635 -95 -2585 1105
rect -2535 -95 -2485 1105
rect -2435 -95 -2385 1105
rect -2335 -95 -2285 1105
rect -2235 -95 -2185 1105
rect -2135 -95 -2085 1105
rect -2035 -95 -1985 1105
rect -1935 -95 -1885 1105
rect -1835 -95 -1785 1105
rect -1735 -95 -1685 1105
rect -1635 -95 -1585 1105
<< nmos >>
rect -2795 1515 -2745 2715
rect -2695 1515 -2645 2715
rect -2620 1515 -2570 2715
rect -2540 1515 -2490 2715
rect -2465 1515 -2415 2715
rect -2385 1515 -2335 2715
rect -2285 1515 -2235 2715
rect -2210 1515 -2160 2715
rect -2135 1515 -2085 2715
rect -2060 1515 -2010 2715
rect -1985 1515 -1935 2715
rect -1885 1515 -1835 2715
rect -2985 -95 -2935 1105
rect -2885 -95 -2835 1105
rect -2785 -95 -2735 1105
rect -2685 -95 -2635 1105
rect -2585 -95 -2535 1105
rect -2485 -95 -2435 1105
rect -2385 -95 -2335 1105
rect -2285 -95 -2235 1105
rect -2185 -95 -2135 1105
rect -2085 -95 -2035 1105
rect -1985 -95 -1935 1105
rect -1885 -95 -1835 1105
rect -1785 -95 -1735 1105
rect -1685 -95 -1635 1105
<< ndiff >>
rect -2845 1515 -2795 2715
rect -2745 1515 -2695 2715
rect -2645 1515 -2620 2715
rect -2570 1515 -2540 2715
rect -2490 1515 -2465 2715
rect -2415 1515 -2385 2715
rect -2335 1515 -2285 2715
rect -2235 1515 -2210 2715
rect -2160 1515 -2135 2715
rect -2085 1515 -2060 2715
rect -2010 1515 -1985 2715
rect -1935 1515 -1885 2715
rect -1835 1515 -1785 2715
rect -3035 1095 -2985 1105
rect -3035 -80 -3025 1095
rect -2995 -80 -2985 1095
rect -3035 -95 -2985 -80
rect -2935 1095 -2885 1105
rect -2935 -80 -2925 1095
rect -2895 -80 -2885 1095
rect -2935 -95 -2885 -80
rect -2835 1095 -2785 1105
rect -2835 -80 -2825 1095
rect -2795 -80 -2785 1095
rect -2835 -95 -2785 -80
rect -2735 1095 -2685 1105
rect -2735 -80 -2725 1095
rect -2695 -80 -2685 1095
rect -2735 -95 -2685 -80
rect -2635 1095 -2585 1105
rect -2635 -80 -2625 1095
rect -2595 -80 -2585 1095
rect -2635 -95 -2585 -80
rect -2535 1095 -2485 1105
rect -2535 -80 -2525 1095
rect -2495 -80 -2485 1095
rect -2535 -95 -2485 -80
rect -2435 1095 -2385 1105
rect -2435 -80 -2425 1095
rect -2395 -80 -2385 1095
rect -2435 -95 -2385 -80
rect -2335 1095 -2285 1105
rect -2335 -80 -2325 1095
rect -2295 -80 -2285 1095
rect -2335 -95 -2285 -80
rect -2235 1095 -2185 1105
rect -2235 -80 -2225 1095
rect -2195 -80 -2185 1095
rect -2235 -95 -2185 -80
rect -2135 1095 -2085 1105
rect -2135 -80 -2125 1095
rect -2095 -80 -2085 1095
rect -2135 -95 -2085 -80
rect -2035 1095 -1985 1105
rect -2035 -80 -2025 1095
rect -1995 -80 -1985 1095
rect -2035 -95 -1985 -80
rect -1935 1095 -1885 1105
rect -1935 -80 -1925 1095
rect -1895 -80 -1885 1095
rect -1935 -95 -1885 -80
rect -1835 1095 -1785 1105
rect -1835 -80 -1825 1095
rect -1795 -80 -1785 1095
rect -1835 -95 -1785 -80
rect -1735 1095 -1685 1105
rect -1735 -80 -1725 1095
rect -1695 -80 -1685 1095
rect -1735 -95 -1685 -80
rect -1635 1095 -1585 1105
rect -1635 -80 -1625 1095
rect -1595 -80 -1585 1095
rect -1635 -95 -1585 -80
<< ndiffc >>
rect -3025 -80 -2995 1095
rect -2925 -80 -2895 1095
rect -2825 -80 -2795 1095
rect -2725 -80 -2695 1095
rect -2625 -80 -2595 1095
rect -2525 -80 -2495 1095
rect -2425 -80 -2395 1095
rect -2325 -80 -2295 1095
rect -2225 -80 -2195 1095
rect -2125 -80 -2095 1095
rect -2025 -80 -1995 1095
rect -1925 -80 -1895 1095
rect -1825 -80 -1795 1095
rect -1725 -80 -1695 1095
rect -1625 -80 -1595 1095
<< poly >>
rect -2795 2715 -2745 2735
rect -2695 2715 -2645 2735
rect -2620 2715 -2570 2735
rect -2540 2715 -2490 2735
rect -2465 2715 -2415 2735
rect -2385 2715 -2335 2735
rect -2285 2715 -2235 2735
rect -2210 2715 -2160 2735
rect -2135 2715 -2085 2735
rect -2060 2715 -2010 2735
rect -1985 2715 -1935 2735
rect -1885 2715 -1835 2735
rect -2795 1495 -2745 1515
rect -2695 1495 -2645 1515
rect -2620 1495 -2570 1515
rect -2540 1495 -2490 1515
rect -2465 1495 -2415 1515
rect -2385 1495 -2335 1515
rect -2285 1495 -2235 1515
rect -2210 1495 -2160 1515
rect -2135 1495 -2085 1515
rect -2060 1495 -2010 1515
rect -1985 1495 -1935 1515
rect -1885 1495 -1835 1515
rect -2985 1105 -2935 1125
rect -2885 1105 -2835 1125
rect -2785 1105 -2735 1125
rect -2685 1105 -2635 1125
rect -2585 1105 -2535 1125
rect -2485 1105 -2435 1125
rect -2385 1105 -2335 1125
rect -2285 1105 -2235 1125
rect -2185 1105 -2135 1125
rect -2085 1105 -2035 1125
rect -1985 1105 -1935 1125
rect -1885 1105 -1835 1125
rect -1785 1105 -1735 1125
rect -1685 1105 -1635 1125
rect -2985 -110 -2935 -95
rect -2885 -110 -2835 -95
rect -2785 -110 -2735 -95
rect -2685 -110 -2635 -95
rect -2585 -110 -2535 -95
rect -2485 -110 -2435 -95
rect -2385 -110 -2335 -95
rect -2285 -110 -2235 -95
rect -2185 -110 -2135 -95
rect -2085 -110 -2035 -95
rect -1985 -110 -1935 -95
rect -1885 -110 -1835 -95
rect -1785 -110 -1735 -95
rect -1685 -110 -1635 -95
<< locali >>
rect -2740 2805 -2700 2820
rect -2740 2755 -2735 2805
rect -2705 2755 -2700 2805
rect -2840 1520 -2800 2715
rect -2740 1525 -2700 2755
rect -1930 2805 -1890 2820
rect -1930 2755 -1925 2805
rect -1895 2755 -1890 2805
rect -2330 1420 -2290 2710
rect -1930 1520 -1890 2755
rect -1830 1520 -1790 2715
rect -3030 1095 -2990 1100
rect -3030 -80 -3025 1095
rect -2995 -80 -2990 1095
rect -3030 -85 -2990 -80
rect -2930 1095 -2890 1100
rect -2930 -80 -2925 1095
rect -2895 -80 -2890 1095
rect -2930 -330 -2890 -80
rect -2830 1095 -2790 1100
rect -2830 -80 -2825 1095
rect -2795 -80 -2790 1095
rect -2830 -85 -2790 -80
rect -2730 1095 -2690 1100
rect -2730 -80 -2725 1095
rect -2695 -80 -2690 1095
rect -2730 -85 -2690 -80
rect -2630 1095 -2590 1100
rect -2630 -80 -2625 1095
rect -2595 -80 -2590 1095
rect -2630 -85 -2590 -80
rect -2530 1095 -2490 1100
rect -2530 -80 -2525 1095
rect -2495 -80 -2490 1095
rect -2530 -85 -2490 -80
rect -2430 1095 -2390 1100
rect -2430 -80 -2425 1095
rect -2395 -80 -2390 1095
rect -2430 -330 -2390 -80
rect -2330 1095 -2290 1100
rect -2330 -80 -2325 1095
rect -2295 -80 -2290 1095
rect -2330 -190 -2290 -80
rect -2230 1095 -2190 1100
rect -2230 -80 -2225 1095
rect -2195 -80 -2190 1095
rect -2230 -330 -2190 -80
rect -2130 1095 -2090 1100
rect -2130 -80 -2125 1095
rect -2095 -80 -2090 1095
rect -2130 -85 -2090 -80
rect -2030 1095 -1990 1100
rect -2030 -80 -2025 1095
rect -1995 -80 -1990 1095
rect -2030 -85 -1990 -80
rect -1930 1095 -1890 1100
rect -1930 -80 -1925 1095
rect -1895 -80 -1890 1095
rect -1930 -85 -1890 -80
rect -1830 1095 -1790 1100
rect -1830 -80 -1825 1095
rect -1795 -80 -1790 1095
rect -1830 -85 -1790 -80
rect -1730 1095 -1690 1100
rect -1730 -80 -1725 1095
rect -1695 -80 -1690 1095
rect -1730 -330 -1690 -80
rect -1630 1095 -1590 1100
rect -1630 -80 -1625 1095
rect -1595 -80 -1590 1095
rect -1630 -85 -1590 -80
<< viali >>
rect -2735 2755 -2705 2805
rect -1925 2755 -1895 2805
<< metal1 >>
rect -2745 2805 -2695 2815
rect -2745 2755 -2735 2805
rect -2705 2800 -2695 2805
rect -1935 2805 -1885 2815
rect -1935 2800 -1925 2805
rect -2705 2760 -1925 2800
rect -2705 2755 -2695 2760
rect -2745 2745 -2695 2755
rect -1935 2755 -1925 2760
rect -1895 2755 -1885 2805
rect -1935 2740 -1885 2755
<< labels >>
flabel locali -2330 -190 -2290 -155 0 FreeSans 800 0 0 0 G
flabel locali -1930 2780 -1890 2810 0 FreeSans 400 0 0 0 VDD
flabel locali -2740 2785 -2700 2815 0 FreeSans 400 0 0 0 VDD
<< end >>
