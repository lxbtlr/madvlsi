magic
tech sky130A
timestamp 1696022310
<< isosubstrate >>
rect -60 862 -4 902
<< nwell >>
rect -210 1040 65 1425
<< locali >>
rect 23 1270 65 1271
rect -30 1250 65 1270
rect -30 1160 -10 1250
rect 35 980 65 1000
rect -199 864 -160 884
rect 35 840 55 980
rect -105 820 55 840
<< metal1 >>
rect 10 1390 65 1425
rect 10 1164 55 1390
rect -204 1069 -195 1164
rect -16 1069 55 1164
rect -15 999 20 1000
rect -204 904 -195 999
rect -16 904 20 999
rect -15 430 20 904
rect -15 350 65 430
use inverte  inverte_0
timestamp 1694482630
transform 1 0 -95 0 1 869
box -110 -30 110 315
use mp2  mp2_0
timestamp 1696021598
transform 1 0 -635 0 1 -75
box 695 295 1115 1500
use mp2  mp2_1
timestamp 1696021598
transform 1 0 -215 0 1 -75
box 695 295 1115 1500
use mp2  mp2_2
timestamp 1696021598
transform 1 0 205 0 1 -75
box 695 295 1115 1500
use mp2  mp2_3
timestamp 1696021598
transform 1 0 625 0 1 -75
box 695 295 1115 1500
<< labels >>
rlabel space 60 845 60 845 7 CLK
port 10 w
rlabel metal1 -204 1112 -204 1112 1 VP
port 6 n
rlabel metal1 -204 949 -204 949 1 VN
port 5 n
rlabel locali -199 875 -199 875 3 D
port 1 e
rlabel space 1740 990 1740 990 3 Q
port 9 e
rlabel space 1740 1255 1740 1255 3 Q_NOT
port 8 e
<< end >>
