* NGSPICE file created from bias_generator.ext - technology: sky130A


* Top level circuit bias_generator

X0 a_n6090_7100# a_n6090_7100# a_n6430_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=6 ps=25 w=12 l=0.5
X1 w_n6530_3120# w_n6530_3120# a_n6230_300# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X2 a_n6030_530# a_n6230_300# a_n6230_300# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X3 a_n4640_8480# a_n5740_8350# a_n5930_11100# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=1.8 pd=12.3 as=3 ps=12.5 w=12 l=0.5
X4 a_n4330_8480# a_n5740_8350# a_n4480_8480# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=1.8 pd=12.3 as=1.5 ps=12.2 w=12 l=0.5
X5 a_n6430_530# a_n5740_8350# a_n4170_8480# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=1.5 ps=12.2 w=12 l=0.5
X6 a_n5930_500# a_n5930_500# a_n5930_500# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=48 ps=200 w=12 l=0.5
X7 a_n5930_11100# a_n5930_11100# a_n6030_11240# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X8 a_n4830_11240# a_n5930_11100# a_n6030_11240# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X9 a_n6430_530# a_n5930_500# a_n6030_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X10 a_n5930_11100# a_n5930_11100# a_n5930_11100# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=48 ps=200 w=12 l=0.5
X11 a_n4990_8480# a_n5740_8350# a_n5140_8480# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X12 a_n6210_6050# a_n6090_7100# a_n6430_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=6 ps=25 w=12 l=0.5
X13 a_n6230_300# w_n6530_3120# w_n6530_3120# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3.6 pd=12.6 as=6 ps=25 w=12 l=0.5
X14 a_n6430_530# a_n6430_530# a_n6230_300# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X15 a_n5140_8480# a_n5740_8350# a_n5290_8480# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X16 a_n6430_530# a_n6090_7100# a_n6210_6050# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3.3 ps=12.6 w=12 l=0.5
X17 a_n6230_11240# a_n5740_8350# a_n6430_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X18 w_n6530_3120# a_n6210_6050# a_n6230_300# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3.6 ps=12.6 w=12 l=0.5
X19 a_n5930_11100# a_n5930_11100# a_n5930_11100# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X20 a_n6030_530# a_n5930_500# a_n5930_500# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X21 a_n6030_11240# a_n5930_11100# a_n4830_11240# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X22 a_n5930_500# a_n5930_500# a_n6030_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X23 a_n6030_11240# a_n5930_11100# a_n5930_11100# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X24 a_n4480_8480# a_n5740_8350# a_n4640_8480# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.8 ps=12.3 w=12 l=0.5
X25 a_n4640_3290# a_n6210_6050# a_n5930_500# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=1.8 pd=12.3 as=3 ps=12.5 w=12 l=0.5
X26 a_n4170_8480# a_n5740_8350# a_n4330_8480# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.8 ps=12.3 w=12 l=0.5
X27 a_n6430_530# a_n6090_7100# a_n6090_7100# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=6 ps=25 w=12 l=0.5
X28 a_n4330_3290# a_n6210_6050# a_n4480_3290# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=1.8 pd=12.3 as=1.5 ps=12.2 w=12 l=0.5
X29 a_n5930_500# a_n5930_500# a_n5930_500# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X30 w_n6530_3120# a_n6210_6050# a_n4170_3290# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=1.5 ps=12.2 w=12 l=0.5
X31 a_n5440_8480# a_n5740_8350# a_n6430_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=3 ps=12.5 w=12 l=0.5
X32 a_n5290_8480# a_n5740_8350# a_n5440_8480# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X33 a_n6230_300# a_n6430_530# a_n6430_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X34 a_n5930_11100# a_n5930_11100# a_n5930_11100# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X35 a_n6230_11240# a_n6430_530# a_n6430_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X36 a_n5140_3290# a_n6210_6050# a_n5290_3290# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X37 a_n4990_3290# a_n6210_6050# a_n5140_3290# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X38 a_n5930_11100# a_n5930_11100# a_n6030_11240# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X39 a_n5930_500# a_n5930_500# a_n5930_500# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X40 a_n6230_11240# a_n6230_11240# a_n6030_11240# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X41 a_n5930_500# a_n5930_500# a_n5930_500# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X42 a_n5930_11100# a_n5740_8350# a_n4990_8480# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=1.5 ps=12.2 w=12 l=0.5
X43 a_n6230_300# a_n6210_6050# w_n6530_3120# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X44 a_n6230_300# a_n6230_300# a_n6030_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X45 a_n6230_11240# w_n6530_3120# w_n6530_3120# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X46 a_n4480_3290# a_n6210_6050# a_n4640_3290# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.8 ps=12.3 w=12 l=0.5
X47 a_n5930_11100# a_n5930_11100# a_n5930_11100# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X48 a_n4170_3290# a_n6210_6050# a_n4330_3290# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.8 ps=12.3 w=12 l=0.5
X49 a_n5930_11100# a_n5930_11100# a_n5930_11100# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X50 w_n6530_3120# w_n6530_3120# a_n6230_11240# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X51 a_n5930_500# a_n5930_500# a_n5930_500# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X52 a_n5290_3290# a_n6210_6050# a_n5440_3290# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X53 a_n6030_530# a_n5930_500# a_n6430_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X54 a_n6430_530# a_n6430_530# a_n6230_11240# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=6 pd=25 as=3 ps=12.5 w=12 l=0.5
X55 a_n5440_3290# a_n6210_6050# w_n6530_3120# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=3 ps=12.5 w=12 l=0.5
X56 a_n6030_11240# a_n6230_11240# a_n6230_11240# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X57 a_n6030_11240# a_n5930_11100# a_n5930_11100# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X58 a_n6210_6050# a_n6210_6050# w_n6530_3120# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=6 pd=25 as=6.6 ps=25.1 w=12 l=0.5
X59 a_n5930_11100# a_n5930_11100# a_n5930_11100# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X60 a_n5930_500# a_n6210_6050# a_n4990_3290# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=3 pd=12.5 as=1.5 ps=12.2 w=12 l=0.5
X61 a_n5930_500# a_n5930_500# a_n6030_530# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X62 a_n5930_500# a_n5930_500# a_n5930_500# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=0 ps=0 w=12 l=0.5
X63 a_n6430_530# a_n5740_8350# a_n6230_11240# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X64 a_n6030_530# a_n5930_500# a_n5930_500# a_n6430_530# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.5
X65 w_n6530_3120# a_n6210_6050# a_n6210_6050# w_n6530_3120# sky130_fd_pr__pfet_01v8 ad=6.6 pd=25.1 as=6 ps=25 w=12 l=0.5
.end

