magic
tech sky130A
timestamp 1697739069
<< nwell >>
rect -3255 5530 -1525 7075
rect -3265 1560 -1535 3375
<< nmos >>
rect -2970 4240 -2920 5440
rect -2870 4240 -2820 5440
rect -2770 4240 -2720 5440
rect -2695 4240 -2645 5440
rect -2620 4240 -2570 5440
rect -2545 4240 -2495 5440
rect -2470 4240 -2420 5440
rect -2370 4240 -2320 5440
rect -2290 4240 -2240 5440
rect -2215 4240 -2165 5440
rect -2135 4240 -2085 5440
rect -2060 4240 -2010 5440
rect -1960 4240 -1910 5440
rect -1860 4240 -1810 5440
rect -3030 4055 -1830 4105
rect -3030 3855 -1830 3905
rect -3030 3750 -1830 3800
rect -3030 3550 -1830 3600
rect -3165 265 -3115 1465
rect -3065 265 -3015 1465
rect -2965 265 -2915 1465
rect -2865 265 -2815 1465
rect -2765 265 -2715 1465
rect -2665 265 -2615 1465
rect -2565 265 -2515 1465
rect -2465 265 -2415 1465
rect -2365 265 -2315 1465
rect -2265 265 -2215 1465
rect -2165 265 -2115 1465
rect -2065 265 -2015 1465
rect -1965 265 -1915 1465
rect -1865 265 -1815 1465
rect -1765 265 -1715 1465
rect -1665 265 -1615 1465
<< pmos >>
rect -3165 5620 -3115 6820
rect -3065 5620 -3015 6820
rect -2965 5620 -2915 6820
rect -2865 5620 -2815 6820
rect -2765 5620 -2715 6820
rect -2665 5620 -2615 6820
rect -2565 5620 -2515 6820
rect -2465 5620 -2415 6820
rect -2365 5620 -2315 6820
rect -2265 5620 -2215 6820
rect -2165 5620 -2115 6820
rect -2065 5620 -2015 6820
rect -1965 5620 -1915 6820
rect -1865 5620 -1815 6820
rect -1765 5620 -1715 6820
rect -1665 5620 -1615 6820
rect -3030 3240 -1830 3290
rect -3030 3025 -1830 3075
rect -2980 1645 -2930 2845
rect -2870 1645 -2820 2845
rect -2770 1645 -2720 2845
rect -2695 1645 -2645 2845
rect -2620 1645 -2570 2845
rect -2545 1645 -2495 2845
rect -2470 1645 -2420 2845
rect -2370 1645 -2320 2845
rect -2290 1645 -2240 2845
rect -2215 1645 -2165 2845
rect -2135 1645 -2085 2845
rect -2060 1645 -2010 2845
rect -1960 1645 -1910 2845
rect -1860 1645 -1810 2845
<< ndiff >>
rect -3020 5425 -2970 5440
rect -3020 4250 -3010 5425
rect -2980 4250 -2970 5425
rect -3020 4240 -2970 4250
rect -2920 5425 -2870 5440
rect -2920 4250 -2910 5425
rect -2880 4250 -2870 5425
rect -2920 4240 -2870 4250
rect -2820 5425 -2770 5440
rect -2820 4250 -2810 5425
rect -2780 4250 -2770 5425
rect -2820 4240 -2770 4250
rect -2720 4240 -2695 5440
rect -2645 4240 -2620 5440
rect -2570 4240 -2545 5440
rect -2495 4240 -2470 5440
rect -2420 5425 -2370 5440
rect -2420 4250 -2410 5425
rect -2380 4250 -2370 5425
rect -2420 4240 -2370 4250
rect -2320 4240 -2290 5440
rect -2240 4240 -2215 5440
rect -2165 4240 -2135 5440
rect -2085 4240 -2060 5440
rect -2010 5425 -1960 5440
rect -2010 4250 -2000 5425
rect -1970 4250 -1960 5425
rect -2010 4240 -1960 4250
rect -1910 5425 -1860 5440
rect -1910 4250 -1900 5425
rect -1870 4250 -1860 5425
rect -1910 4240 -1860 4250
rect -1810 5425 -1760 5440
rect -1810 4250 -1800 5425
rect -1770 4250 -1760 5425
rect -1810 4240 -1760 4250
rect -3030 4145 -1830 4155
rect -3030 4115 -3020 4145
rect -1845 4115 -1830 4145
rect -3030 4105 -1830 4115
rect -3030 4045 -1830 4055
rect -3030 4015 -3020 4045
rect -1845 4015 -1830 4045
rect -3030 4005 -1830 4015
rect -3030 3945 -1830 3955
rect -3030 3915 -3020 3945
rect -1845 3915 -1830 3945
rect -3030 3905 -1830 3915
rect -3030 3845 -1830 3855
rect -3030 3810 -3020 3845
rect -1845 3810 -1830 3845
rect -3030 3800 -1830 3810
rect -3030 3740 -1830 3750
rect -3030 3710 -3020 3740
rect -1845 3710 -1830 3740
rect -3030 3700 -1830 3710
rect -3030 3640 -1830 3650
rect -3030 3610 -3020 3640
rect -1845 3610 -1830 3640
rect -3030 3600 -1830 3610
rect -3030 3540 -1830 3550
rect -3030 3510 -3020 3540
rect -1845 3510 -1830 3540
rect -3030 3500 -1830 3510
rect -3215 1455 -3165 1465
rect -3215 280 -3205 1455
rect -3175 280 -3165 1455
rect -3215 265 -3165 280
rect -3115 1455 -3065 1465
rect -3115 280 -3105 1455
rect -3075 280 -3065 1455
rect -3115 265 -3065 280
rect -3015 1455 -2965 1465
rect -3015 280 -3005 1455
rect -2975 280 -2965 1455
rect -3015 265 -2965 280
rect -2915 1455 -2865 1465
rect -2915 280 -2905 1455
rect -2875 280 -2865 1455
rect -2915 265 -2865 280
rect -2815 1455 -2765 1465
rect -2815 280 -2805 1455
rect -2775 280 -2765 1455
rect -2815 265 -2765 280
rect -2715 1455 -2665 1465
rect -2715 280 -2705 1455
rect -2675 280 -2665 1455
rect -2715 265 -2665 280
rect -2615 1455 -2565 1465
rect -2615 280 -2605 1455
rect -2575 280 -2565 1455
rect -2615 265 -2565 280
rect -2515 1455 -2465 1465
rect -2515 280 -2505 1455
rect -2475 280 -2465 1455
rect -2515 265 -2465 280
rect -2415 1455 -2365 1465
rect -2415 280 -2405 1455
rect -2375 280 -2365 1455
rect -2415 265 -2365 280
rect -2315 1455 -2265 1465
rect -2315 280 -2305 1455
rect -2275 280 -2265 1455
rect -2315 265 -2265 280
rect -2215 1455 -2165 1465
rect -2215 280 -2205 1455
rect -2175 280 -2165 1455
rect -2215 265 -2165 280
rect -2115 1455 -2065 1465
rect -2115 280 -2105 1455
rect -2075 280 -2065 1455
rect -2115 265 -2065 280
rect -2015 1455 -1965 1465
rect -2015 280 -2005 1455
rect -1975 280 -1965 1455
rect -2015 265 -1965 280
rect -1915 1455 -1865 1465
rect -1915 280 -1905 1455
rect -1875 280 -1865 1455
rect -1915 265 -1865 280
rect -1815 1455 -1765 1465
rect -1815 280 -1805 1455
rect -1775 280 -1765 1455
rect -1815 265 -1765 280
rect -1715 1455 -1665 1465
rect -1715 280 -1705 1455
rect -1675 280 -1665 1455
rect -1715 265 -1665 280
rect -1615 1455 -1565 1465
rect -1615 280 -1605 1455
rect -1575 280 -1565 1455
rect -1615 265 -1565 280
<< pdiff >>
rect -3215 6805 -3165 6820
rect -3215 5630 -3205 6805
rect -3175 5630 -3165 6805
rect -3215 5620 -3165 5630
rect -3115 6805 -3065 6820
rect -3115 5630 -3105 6805
rect -3075 5630 -3065 6805
rect -3115 5620 -3065 5630
rect -3015 6805 -2965 6820
rect -3015 5630 -3005 6805
rect -2975 5630 -2965 6805
rect -3015 5620 -2965 5630
rect -2915 6805 -2865 6820
rect -2915 5630 -2905 6805
rect -2875 5630 -2865 6805
rect -2915 5620 -2865 5630
rect -2815 6805 -2765 6820
rect -2815 5630 -2805 6805
rect -2775 5630 -2765 6805
rect -2815 5620 -2765 5630
rect -2715 6805 -2665 6820
rect -2715 5630 -2705 6805
rect -2675 5630 -2665 6805
rect -2715 5620 -2665 5630
rect -2615 6805 -2565 6820
rect -2615 5630 -2605 6805
rect -2575 5630 -2565 6805
rect -2615 5620 -2565 5630
rect -2515 6805 -2465 6820
rect -2515 5630 -2505 6805
rect -2475 5630 -2465 6805
rect -2515 5620 -2465 5630
rect -2415 6805 -2365 6820
rect -2415 5630 -2405 6805
rect -2375 5630 -2365 6805
rect -2415 5620 -2365 5630
rect -2315 6805 -2265 6820
rect -2315 5630 -2305 6805
rect -2275 5630 -2265 6805
rect -2315 5620 -2265 5630
rect -2215 6805 -2165 6820
rect -2215 5630 -2205 6805
rect -2175 5630 -2165 6805
rect -2215 5620 -2165 5630
rect -2115 6805 -2065 6820
rect -2115 5630 -2105 6805
rect -2075 5630 -2065 6805
rect -2115 5620 -2065 5630
rect -2015 6805 -1965 6820
rect -2015 5630 -2005 6805
rect -1975 5630 -1965 6805
rect -2015 5620 -1965 5630
rect -1915 6805 -1865 6820
rect -1915 5630 -1905 6805
rect -1875 5630 -1865 6805
rect -1915 5620 -1865 5630
rect -1815 6805 -1765 6820
rect -1815 5630 -1805 6805
rect -1775 5630 -1765 6805
rect -1815 5620 -1765 5630
rect -1715 6805 -1665 6820
rect -1715 5630 -1705 6805
rect -1675 5630 -1665 6805
rect -1715 5620 -1665 5630
rect -1615 6805 -1565 6820
rect -1615 5630 -1605 6805
rect -1575 5630 -1565 6805
rect -1615 5620 -1565 5630
rect -3030 3330 -1830 3340
rect -3030 3300 -3020 3330
rect -1845 3300 -1830 3330
rect -3030 3290 -1830 3300
rect -3030 3230 -1830 3240
rect -3030 3195 -3020 3230
rect -1845 3195 -1830 3230
rect -3030 3185 -1830 3195
rect -3030 3120 -1830 3130
rect -3030 3085 -3020 3120
rect -1845 3085 -1830 3120
rect -3030 3075 -1830 3085
rect -3030 3015 -1830 3025
rect -3030 2985 -3020 3015
rect -1845 2985 -1830 3015
rect -3030 2975 -1830 2985
rect -3030 2835 -2980 2845
rect -3030 1660 -3020 2835
rect -2990 1660 -2980 2835
rect -3030 1645 -2980 1660
rect -2930 2835 -2870 2845
rect -2930 1660 -2920 2835
rect -2880 1660 -2870 2835
rect -2930 1645 -2870 1660
rect -2820 2835 -2770 2845
rect -2820 1660 -2810 2835
rect -2780 1660 -2770 2835
rect -2820 1645 -2770 1660
rect -2720 1645 -2695 2845
rect -2645 1645 -2620 2845
rect -2570 1645 -2545 2845
rect -2495 1645 -2470 2845
rect -2420 2835 -2370 2845
rect -2420 1660 -2410 2835
rect -2380 1660 -2370 2835
rect -2420 1645 -2370 1660
rect -2320 1645 -2290 2845
rect -2240 1645 -2215 2845
rect -2165 1645 -2135 2845
rect -2085 1645 -2060 2845
rect -2010 2835 -1960 2845
rect -2010 1660 -2000 2835
rect -1970 1660 -1960 2835
rect -2010 1645 -1960 1660
rect -1910 2835 -1860 2845
rect -1910 1660 -1900 2835
rect -1870 1660 -1860 2835
rect -1910 1645 -1860 1660
rect -1810 2835 -1760 2845
rect -1810 1660 -1800 2835
rect -1770 1660 -1760 2835
rect -1810 1645 -1760 1660
<< ndiffc >>
rect -3010 4250 -2980 5425
rect -2910 4250 -2880 5425
rect -2810 4250 -2780 5425
rect -2410 4250 -2380 5425
rect -2000 4250 -1970 5425
rect -1900 4250 -1870 5425
rect -1800 4250 -1770 5425
rect -3020 4115 -1845 4145
rect -3020 4015 -1845 4045
rect -3020 3915 -1845 3945
rect -3020 3810 -1845 3845
rect -3020 3710 -1845 3740
rect -3020 3610 -1845 3640
rect -3020 3510 -1845 3540
rect -3205 280 -3175 1455
rect -3105 280 -3075 1455
rect -3005 280 -2975 1455
rect -2905 280 -2875 1455
rect -2805 280 -2775 1455
rect -2705 280 -2675 1455
rect -2605 280 -2575 1455
rect -2505 280 -2475 1455
rect -2405 280 -2375 1455
rect -2305 280 -2275 1455
rect -2205 280 -2175 1455
rect -2105 280 -2075 1455
rect -2005 280 -1975 1455
rect -1905 280 -1875 1455
rect -1805 280 -1775 1455
rect -1705 280 -1675 1455
rect -1605 280 -1575 1455
<< pdiffc >>
rect -3205 5630 -3175 6805
rect -3105 5630 -3075 6805
rect -3005 5630 -2975 6805
rect -2905 5630 -2875 6805
rect -2805 5630 -2775 6805
rect -2705 5630 -2675 6805
rect -2605 5630 -2575 6805
rect -2505 5630 -2475 6805
rect -2405 5630 -2375 6805
rect -2305 5630 -2275 6805
rect -2205 5630 -2175 6805
rect -2105 5630 -2075 6805
rect -2005 5630 -1975 6805
rect -1905 5630 -1875 6805
rect -1805 5630 -1775 6805
rect -1705 5630 -1675 6805
rect -1605 5630 -1575 6805
rect -3020 3300 -1845 3330
rect -3020 3195 -1845 3230
rect -3020 3085 -1845 3120
rect -3020 2985 -1845 3015
rect -3020 1660 -2990 2835
rect -2920 1660 -2880 2835
rect -2810 1660 -2780 2835
rect -2410 1660 -2380 2835
rect -2000 1660 -1970 2835
rect -1900 1660 -1870 2835
rect -1800 1660 -1770 2835
<< psubdiff >>
rect -3070 5420 -3020 5440
rect -3070 4255 -3060 5420
rect -3030 4255 -3020 5420
rect -3070 4240 -3020 4255
rect -1760 5425 -1710 5440
rect -1760 4255 -1750 5425
rect -1720 4255 -1710 5425
rect -1760 4240 -1710 4255
rect -3030 3995 -1830 4005
rect -3030 3965 -3020 3995
rect -1845 3965 -1830 3995
rect -3030 3955 -1830 3965
rect -3030 3690 -1830 3700
rect -3030 3660 -3020 3690
rect -1845 3660 -1830 3690
rect -3030 3650 -1830 3660
rect -2955 80 -1755 95
rect -2955 60 -2940 80
rect -1780 60 -1755 80
rect -2955 45 -1755 60
<< nsubdiff >>
rect -2990 7035 -1790 7050
rect -2990 7005 -2980 7035
rect -1800 7005 -1790 7035
rect -2990 6990 -1790 7005
rect -3030 3175 -1830 3185
rect -3030 3140 -3020 3175
rect -1845 3140 -1830 3175
rect -3030 3130 -1830 3140
rect -3080 2830 -3030 2845
rect -3080 1665 -3070 2830
rect -3040 1665 -3030 2830
rect -3080 1645 -3030 1665
rect -1760 2830 -1710 2845
rect -1760 1665 -1750 2830
rect -1720 1665 -1710 2830
rect -1760 1645 -1710 1665
<< psubdiffcont >>
rect -3060 4255 -3030 5420
rect -1750 4255 -1720 5425
rect -3020 3965 -1845 3995
rect -3020 3660 -1845 3690
rect -2940 60 -1780 80
<< nsubdiffcont >>
rect -2980 7005 -1800 7035
rect -3020 3140 -1845 3175
rect -3070 1665 -3040 2830
rect -1750 1665 -1720 2830
<< poly >>
rect -3115 6925 -3015 6935
rect -3115 6895 -3105 6925
rect -3075 6895 -3015 6925
rect -3115 6885 -3015 6895
rect -3165 6820 -3115 6835
rect -3065 6820 -3015 6885
rect -1765 6925 -1665 6935
rect -1765 6895 -1705 6925
rect -1675 6895 -1665 6925
rect -1765 6885 -1665 6895
rect -2965 6820 -2915 6835
rect -2865 6820 -2815 6835
rect -2765 6820 -2715 6835
rect -2665 6820 -2615 6835
rect -2565 6820 -2515 6835
rect -2465 6820 -2415 6835
rect -2365 6820 -2315 6835
rect -2265 6820 -2215 6835
rect -2165 6820 -2115 6835
rect -2065 6820 -2015 6835
rect -1965 6820 -1915 6835
rect -1865 6820 -1815 6835
rect -1765 6820 -1715 6885
rect -1665 6820 -1615 6835
rect -3165 5600 -3115 5620
rect -3215 5590 -3115 5600
rect -3215 5560 -3205 5590
rect -3175 5560 -3115 5590
rect -3215 5550 -3115 5560
rect -3065 5590 -3015 5620
rect -3065 5560 -3055 5590
rect -3025 5560 -3015 5590
rect -3065 5550 -3015 5560
rect -2965 5590 -2915 5620
rect -2965 5560 -2955 5590
rect -2925 5560 -2915 5590
rect -2965 5550 -2915 5560
rect -2865 5590 -2815 5620
rect -2865 5560 -2855 5590
rect -2825 5560 -2815 5590
rect -2865 5550 -2815 5560
rect -2765 5590 -2715 5620
rect -2765 5560 -2755 5590
rect -2725 5560 -2715 5590
rect -2765 5550 -2715 5560
rect -2665 5590 -2615 5620
rect -2665 5560 -2655 5590
rect -2625 5560 -2615 5590
rect -2665 5550 -2615 5560
rect -2565 5590 -2515 5620
rect -2565 5560 -2555 5590
rect -2525 5560 -2515 5590
rect -2565 5550 -2515 5560
rect -2465 5590 -2415 5620
rect -2465 5560 -2455 5590
rect -2425 5560 -2415 5590
rect -2465 5550 -2415 5560
rect -2365 5590 -2315 5620
rect -2365 5560 -2355 5590
rect -2325 5560 -2315 5590
rect -2365 5550 -2315 5560
rect -2265 5590 -2215 5620
rect -2265 5560 -2255 5590
rect -2225 5560 -2215 5590
rect -2265 5550 -2215 5560
rect -2165 5590 -2115 5620
rect -2165 5560 -2155 5590
rect -2125 5560 -2115 5590
rect -2165 5550 -2115 5560
rect -2065 5590 -2015 5620
rect -2065 5560 -2055 5590
rect -2025 5560 -2015 5590
rect -2065 5550 -2015 5560
rect -1965 5590 -1915 5620
rect -1965 5560 -1955 5590
rect -1925 5560 -1915 5590
rect -1965 5550 -1915 5560
rect -1865 5590 -1815 5620
rect -1865 5560 -1855 5590
rect -1825 5560 -1815 5590
rect -1865 5550 -1815 5560
rect -1765 5590 -1715 5620
rect -1765 5560 -1755 5590
rect -1725 5560 -1715 5590
rect -1765 5550 -1715 5560
rect -1665 5600 -1615 5620
rect -1665 5590 -1565 5600
rect -1665 5560 -1605 5590
rect -1575 5560 -1565 5590
rect -1665 5550 -1565 5560
rect -2970 5440 -2920 5455
rect -2870 5440 -2820 5460
rect -2770 5440 -2720 5460
rect -2695 5440 -2645 5460
rect -2620 5440 -2570 5460
rect -2545 5440 -2495 5460
rect -2470 5440 -2420 5460
rect -2370 5440 -2320 5460
rect -2290 5440 -2240 5460
rect -2215 5440 -2165 5460
rect -2135 5440 -2085 5460
rect -2060 5440 -2010 5460
rect -1960 5440 -1910 5460
rect -1860 5440 -1810 5455
rect -2970 4220 -2920 4240
rect -3020 4210 -2920 4220
rect -3020 4180 -3010 4210
rect -2980 4180 -2920 4210
rect -3020 4170 -2920 4180
rect -2870 4220 -2820 4240
rect -2770 4220 -2720 4240
rect -2695 4220 -2645 4240
rect -2620 4220 -2570 4240
rect -2545 4220 -2495 4240
rect -2470 4220 -2420 4240
rect -2370 4220 -2320 4240
rect -2290 4220 -2240 4240
rect -2215 4220 -2165 4240
rect -2135 4220 -2085 4240
rect -2060 4220 -2010 4240
rect -1960 4220 -1910 4240
rect -2870 4210 -1910 4220
rect -2870 4180 -2410 4210
rect -2380 4180 -1950 4210
rect -1920 4180 -1910 4210
rect -2870 4175 -1910 4180
rect -2420 4170 -2370 4175
rect -1960 4170 -1910 4175
rect -1860 4220 -1810 4240
rect -1860 4210 -1760 4220
rect -1860 4180 -1800 4210
rect -1770 4180 -1760 4210
rect -1860 4170 -1760 4180
rect -3045 4055 -3030 4105
rect -1830 4095 -1760 4105
rect -1830 4065 -1800 4095
rect -1770 4065 -1760 4095
rect -1830 4055 -1760 4065
rect -1810 3905 -1760 4055
rect -3045 3855 -3030 3905
rect -1830 3855 -1760 3905
rect -1810 3800 -1760 3855
rect -3045 3750 -3030 3800
rect -1830 3750 -1760 3800
rect -1810 3600 -1760 3750
rect -3045 3550 -3030 3600
rect -1830 3590 -1760 3600
rect -1830 3560 -1800 3590
rect -1770 3560 -1760 3590
rect -1830 3550 -1760 3560
rect -3105 3280 -3030 3290
rect -3105 3250 -3095 3280
rect -3065 3250 -3030 3280
rect -3105 3240 -3030 3250
rect -1830 3240 -1810 3290
rect -3105 3065 -3030 3075
rect -3105 3035 -3095 3065
rect -3065 3035 -3030 3065
rect -3105 3025 -3030 3035
rect -1830 3025 -1810 3075
rect -3030 2905 -2930 2915
rect -3030 2875 -3020 2905
rect -2990 2875 -2930 2905
rect -2695 2905 -2645 2915
rect -2695 2890 -2685 2905
rect -3030 2865 -2930 2875
rect -2980 2845 -2930 2865
rect -2870 2875 -2685 2890
rect -2655 2890 -2645 2905
rect -1860 2905 -1760 2915
rect -2655 2875 -1910 2890
rect -2870 2865 -1910 2875
rect -2870 2845 -2820 2865
rect -2770 2845 -2720 2865
rect -2695 2845 -2645 2865
rect -2620 2845 -2570 2865
rect -2545 2845 -2495 2865
rect -2470 2845 -2420 2865
rect -2370 2845 -2320 2865
rect -2290 2845 -2240 2865
rect -2215 2845 -2165 2865
rect -2135 2845 -2085 2865
rect -2060 2845 -2010 2865
rect -1960 2845 -1910 2865
rect -1860 2875 -1800 2905
rect -1770 2875 -1760 2905
rect -1860 2865 -1760 2875
rect -1860 2845 -1810 2865
rect -2980 1630 -2930 1645
rect -2870 1625 -2820 1645
rect -2770 1625 -2720 1645
rect -2695 1625 -2645 1645
rect -2620 1625 -2570 1645
rect -2545 1625 -2495 1645
rect -2470 1625 -2420 1645
rect -2370 1625 -2320 1645
rect -2290 1625 -2240 1645
rect -2215 1625 -2165 1645
rect -2135 1625 -2085 1645
rect -2060 1625 -2010 1645
rect -1960 1625 -1910 1645
rect -1860 1630 -1810 1645
rect -3215 1525 -3115 1535
rect -3215 1495 -3205 1525
rect -3175 1495 -3115 1525
rect -3215 1485 -3115 1495
rect -3165 1465 -3115 1485
rect -3065 1525 -3015 1535
rect -3065 1495 -3055 1525
rect -3025 1495 -3015 1525
rect -3065 1465 -3015 1495
rect -2965 1525 -2915 1535
rect -2965 1495 -2955 1525
rect -2925 1495 -2915 1525
rect -2965 1465 -2915 1495
rect -2865 1525 -2815 1535
rect -2865 1495 -2855 1525
rect -2825 1495 -2815 1525
rect -2865 1465 -2815 1495
rect -2765 1525 -2715 1535
rect -2765 1495 -2755 1525
rect -2725 1495 -2715 1525
rect -2765 1465 -2715 1495
rect -2665 1525 -2615 1535
rect -2665 1495 -2655 1525
rect -2625 1495 -2615 1525
rect -2665 1465 -2615 1495
rect -2565 1525 -2515 1535
rect -2565 1495 -2555 1525
rect -2525 1495 -2515 1525
rect -2565 1465 -2515 1495
rect -2465 1525 -2415 1535
rect -2465 1495 -2455 1525
rect -2425 1495 -2415 1525
rect -2465 1465 -2415 1495
rect -2365 1525 -2315 1535
rect -2365 1495 -2355 1525
rect -2325 1495 -2315 1525
rect -2365 1465 -2315 1495
rect -2265 1525 -2215 1535
rect -2265 1495 -2255 1525
rect -2225 1495 -2215 1525
rect -2265 1465 -2215 1495
rect -2165 1525 -2115 1535
rect -2165 1495 -2155 1525
rect -2125 1495 -2115 1525
rect -2165 1465 -2115 1495
rect -2065 1525 -2015 1535
rect -2065 1495 -2055 1525
rect -2025 1495 -2015 1525
rect -2065 1465 -2015 1495
rect -1965 1525 -1915 1535
rect -1965 1495 -1955 1525
rect -1925 1495 -1915 1525
rect -1965 1465 -1915 1495
rect -1865 1525 -1815 1535
rect -1865 1495 -1855 1525
rect -1825 1495 -1815 1525
rect -1865 1465 -1815 1495
rect -1765 1525 -1715 1535
rect -1765 1495 -1755 1525
rect -1725 1495 -1715 1525
rect -1765 1465 -1715 1495
rect -1665 1525 -1565 1535
rect -1665 1495 -1605 1525
rect -1575 1495 -1565 1525
rect -1665 1485 -1565 1495
rect -1665 1465 -1615 1485
rect -3165 250 -3115 265
rect -3065 200 -3015 265
rect -2965 250 -2915 265
rect -2865 250 -2815 265
rect -2765 250 -2715 265
rect -2665 250 -2615 265
rect -2565 250 -2515 265
rect -2465 250 -2415 265
rect -2365 250 -2315 265
rect -2265 250 -2215 265
rect -2165 250 -2115 265
rect -2065 250 -2015 265
rect -1965 250 -1915 265
rect -1865 250 -1815 265
rect -3115 190 -3015 200
rect -3115 160 -3105 190
rect -3075 160 -3015 190
rect -3115 150 -3015 160
rect -1765 200 -1715 265
rect -1665 250 -1615 265
rect -1765 190 -1665 200
rect -1765 160 -1705 190
rect -1675 160 -1665 190
rect -1765 150 -1665 160
<< polycont >>
rect -3105 6895 -3075 6925
rect -1705 6895 -1675 6925
rect -3205 5560 -3175 5590
rect -3055 5560 -3025 5590
rect -2955 5560 -2925 5590
rect -2855 5560 -2825 5590
rect -2755 5560 -2725 5590
rect -2655 5560 -2625 5590
rect -2555 5560 -2525 5590
rect -2455 5560 -2425 5590
rect -2355 5560 -2325 5590
rect -2255 5560 -2225 5590
rect -2155 5560 -2125 5590
rect -2055 5560 -2025 5590
rect -1955 5560 -1925 5590
rect -1855 5560 -1825 5590
rect -1755 5560 -1725 5590
rect -1605 5560 -1575 5590
rect -3010 4180 -2980 4210
rect -2410 4180 -2380 4210
rect -1950 4180 -1920 4210
rect -1800 4180 -1770 4210
rect -1800 4065 -1770 4095
rect -1800 3560 -1770 3590
rect -3095 3250 -3065 3280
rect -3095 3035 -3065 3065
rect -3020 2875 -2990 2905
rect -2685 2875 -2655 2905
rect -1800 2875 -1770 2905
rect -3205 1495 -3175 1525
rect -3055 1495 -3025 1525
rect -2955 1495 -2925 1525
rect -2855 1495 -2825 1525
rect -2755 1495 -2725 1525
rect -2655 1495 -2625 1525
rect -2555 1495 -2525 1525
rect -2455 1495 -2425 1525
rect -2355 1495 -2325 1525
rect -2255 1495 -2225 1525
rect -2155 1495 -2125 1525
rect -2055 1495 -2025 1525
rect -1955 1495 -1925 1525
rect -1855 1495 -1825 1525
rect -1755 1495 -1725 1525
rect -1605 1495 -1575 1525
rect -3105 160 -3075 190
rect -1705 160 -1675 190
<< locali >>
rect -2990 7035 -1790 7045
rect -2990 7005 -2980 7035
rect -1800 7005 -1790 7035
rect -2990 6995 -1790 7005
rect -3110 6935 -1670 6965
rect -3115 6925 -1665 6935
rect -3115 6895 -3105 6925
rect -3075 6895 -3065 6925
rect -3115 6885 -3065 6895
rect -1715 6895 -1705 6925
rect -1675 6895 -1665 6925
rect -1715 6885 -1665 6895
rect -3210 6805 -3170 6820
rect -3210 5630 -3205 6805
rect -3175 5630 -3170 6805
rect -3210 5620 -3170 5630
rect -3110 6805 -3070 6885
rect -3010 6845 -1770 6885
rect -3010 6820 -2970 6845
rect -2510 6820 -2470 6845
rect -2310 6820 -2270 6845
rect -1810 6820 -1770 6845
rect -3110 5630 -3105 6805
rect -3075 5630 -3070 6805
rect -3110 5625 -3070 5630
rect -3205 5600 -3175 5620
rect -3105 5600 -3070 5625
rect -3015 6805 -2965 6820
rect -3015 5630 -3005 6805
rect -2975 5630 -2965 6805
rect -3015 5620 -2965 5630
rect -2915 6805 -2865 6820
rect -2915 5630 -2905 6805
rect -2875 5630 -2865 6805
rect -2915 5620 -2865 5630
rect -2815 6805 -2765 6820
rect -2815 5630 -2805 6805
rect -2775 5630 -2765 6805
rect -2815 5620 -2765 5630
rect -2715 6805 -2665 6820
rect -2715 5630 -2705 6805
rect -2675 5630 -2665 6805
rect -2715 5620 -2665 5630
rect -2615 6805 -2565 6820
rect -2615 5630 -2605 6805
rect -2575 5630 -2565 6805
rect -2615 5620 -2565 5630
rect -2515 6805 -2465 6820
rect -2515 5630 -2505 6805
rect -2475 5630 -2465 6805
rect -2515 5620 -2465 5630
rect -2415 6805 -2365 6820
rect -2415 5630 -2405 6805
rect -2375 5630 -2365 6805
rect -2415 5620 -2365 5630
rect -2315 6805 -2265 6820
rect -2315 5630 -2305 6805
rect -2275 5630 -2265 6805
rect -2315 5620 -2265 5630
rect -2215 6805 -2165 6820
rect -2215 5630 -2205 6805
rect -2175 5630 -2165 6805
rect -2215 5620 -2165 5630
rect -2115 6805 -2065 6820
rect -2115 5630 -2105 6805
rect -2075 5630 -2065 6805
rect -2115 5620 -2065 5630
rect -2015 6805 -1965 6820
rect -2015 5630 -2005 6805
rect -1975 5630 -1965 6805
rect -2015 5620 -1965 5630
rect -1915 6805 -1865 6820
rect -1915 5630 -1905 6805
rect -1875 5630 -1865 6805
rect -1915 5620 -1865 5630
rect -1815 6805 -1765 6820
rect -1815 5630 -1805 6805
rect -1775 5630 -1765 6805
rect -1815 5620 -1765 5630
rect -1710 6805 -1670 6885
rect -1710 5630 -1705 6805
rect -1675 5630 -1670 6805
rect -1710 5625 -1670 5630
rect -1610 6805 -1570 6820
rect -1610 5630 -1605 6805
rect -1575 5630 -1570 6805
rect -2905 5600 -2875 5620
rect -2805 5600 -2775 5620
rect -2705 5600 -2675 5620
rect -2605 5600 -2575 5620
rect -2205 5600 -2175 5620
rect -2105 5600 -2075 5620
rect -2005 5600 -1975 5620
rect -1905 5600 -1875 5620
rect -1710 5600 -1675 5625
rect -1610 5620 -1570 5630
rect -1605 5600 -1575 5620
rect -3215 5590 -3165 5600
rect -3215 5560 -3205 5590
rect -3175 5560 -3165 5590
rect -3215 5550 -3165 5560
rect -3105 5590 -3015 5600
rect -3105 5560 -3055 5590
rect -3025 5560 -3015 5590
rect -3105 5550 -3015 5560
rect -2965 5590 -2515 5600
rect -2965 5560 -2955 5590
rect -2925 5565 -2855 5590
rect -2925 5560 -2915 5565
rect -2965 5550 -2915 5560
rect -2865 5560 -2855 5565
rect -2825 5565 -2755 5590
rect -2825 5560 -2815 5565
rect -2865 5550 -2815 5560
rect -2765 5560 -2755 5565
rect -2725 5565 -2655 5590
rect -2725 5560 -2715 5565
rect -2765 5550 -2715 5560
rect -2665 5560 -2655 5565
rect -2625 5565 -2555 5590
rect -2625 5560 -2615 5565
rect -2665 5550 -2615 5560
rect -2565 5560 -2555 5565
rect -2525 5585 -2515 5590
rect -2465 5590 -2415 5600
rect -2465 5585 -2455 5590
rect -2525 5560 -2455 5585
rect -2425 5585 -2415 5590
rect -2365 5590 -2315 5600
rect -2365 5585 -2355 5590
rect -2425 5560 -2355 5585
rect -2325 5585 -2315 5590
rect -2265 5590 -1815 5600
rect -2265 5585 -2255 5590
rect -2325 5560 -2255 5585
rect -2225 5565 -2155 5590
rect -2225 5560 -2215 5565
rect -2565 5550 -2215 5560
rect -2165 5560 -2155 5565
rect -2125 5565 -2055 5590
rect -2125 5560 -2115 5565
rect -2165 5550 -2115 5560
rect -2065 5560 -2055 5565
rect -2025 5565 -1955 5590
rect -2025 5560 -2015 5565
rect -2065 5550 -2015 5560
rect -1965 5560 -1955 5565
rect -1925 5565 -1855 5590
rect -1925 5560 -1915 5565
rect -1965 5550 -1915 5560
rect -1865 5560 -1855 5565
rect -1825 5560 -1815 5590
rect -1865 5550 -1815 5560
rect -1765 5590 -1675 5600
rect -1765 5560 -1755 5590
rect -1725 5560 -1675 5590
rect -1765 5550 -1675 5560
rect -1615 5590 -1565 5600
rect -1615 5560 -1605 5590
rect -1575 5560 -1565 5590
rect -1615 5550 -1565 5560
rect -3105 5510 -3070 5550
rect -3105 5470 -2875 5510
rect -3070 5425 -2975 5440
rect -3070 5420 -3010 5425
rect -3070 4255 -3060 5420
rect -3030 4255 -3010 5420
rect -3070 4250 -3010 4255
rect -2980 4250 -2975 5425
rect -3070 4240 -2975 4250
rect -2915 5425 -2875 5470
rect -2915 4250 -2910 5425
rect -2880 4250 -2875 5425
rect -2915 4240 -2875 4250
rect -2815 5425 -2775 5435
rect -2815 4250 -2810 5425
rect -2780 4250 -2775 5425
rect -2815 4240 -2775 4250
rect -2415 5425 -2375 5550
rect -1710 5510 -1675 5550
rect -1905 5470 -1675 5510
rect -2415 4250 -2410 5425
rect -2380 4250 -2375 5425
rect -2415 4240 -2375 4250
rect -2005 5425 -1965 5435
rect -2005 4250 -2000 5425
rect -1970 4250 -1965 5425
rect -2005 4240 -1965 4250
rect -1905 5425 -1865 5470
rect -1905 4250 -1900 5425
rect -1870 4250 -1865 5425
rect -1905 4240 -1865 4250
rect -1805 5425 -1705 5440
rect -1805 4250 -1800 5425
rect -1770 4255 -1750 5425
rect -1720 4255 -1705 5425
rect -1770 4250 -1705 4255
rect -1805 4240 -1705 4250
rect -3010 4220 -2980 4240
rect -1800 4220 -1770 4240
rect -3020 4210 -2970 4220
rect -3020 4180 -3010 4210
rect -2980 4180 -2970 4210
rect -3020 4170 -2970 4180
rect -2420 4210 -2370 4220
rect -2420 4180 -2410 4210
rect -2380 4180 -2370 4210
rect -2420 4170 -2370 4180
rect -1960 4210 -1910 4220
rect -1960 4180 -1950 4210
rect -1920 4180 -1910 4210
rect -1960 4170 -1910 4180
rect -1810 4210 -1760 4220
rect -1810 4180 -1800 4210
rect -1770 4180 -1760 4210
rect -1810 4170 -1760 4180
rect -3030 4145 -1840 4150
rect -3030 4115 -3020 4145
rect -1845 4115 -1780 4145
rect -3030 4110 -1840 4115
rect -1810 4105 -1780 4115
rect -1810 4095 -1760 4105
rect -1810 4065 -1800 4095
rect -1770 4065 -1760 4095
rect -1810 4055 -1760 4065
rect -3030 4045 -1835 4050
rect -3030 4015 -3020 4045
rect -1845 4015 -1835 4045
rect -3030 3995 -1835 4015
rect -3030 3965 -3020 3995
rect -1845 3965 -1835 3995
rect -3030 3945 -1835 3965
rect -3030 3915 -3020 3945
rect -1845 3915 -1835 3945
rect -3030 3910 -1835 3915
rect -3095 3845 -1835 3850
rect -3095 3810 -3020 3845
rect -1845 3810 -1835 3845
rect -3095 3805 -1835 3810
rect -3095 3335 -3050 3805
rect -3030 3740 -1835 3745
rect -3030 3710 -3020 3740
rect -1845 3710 -1835 3740
rect -3030 3690 -1835 3710
rect -3030 3660 -3020 3690
rect -1845 3660 -1835 3690
rect -3030 3640 -1835 3660
rect -3030 3610 -3020 3640
rect -1845 3610 -1835 3640
rect -3030 3605 -1835 3610
rect -1810 3590 -1760 3600
rect -1810 3560 -1800 3590
rect -1770 3560 -1760 3590
rect -1810 3550 -1760 3560
rect -3030 3540 -1840 3545
rect -1810 3540 -1780 3550
rect -3030 3510 -3020 3540
rect -1845 3510 -1780 3540
rect -3030 3505 -1840 3510
rect -3095 3330 -1835 3335
rect -3095 3300 -3020 3330
rect -1845 3300 -1835 3330
rect -3095 3295 -1835 3300
rect -3095 3290 -3055 3295
rect -3105 3280 -3055 3290
rect -3105 3250 -3095 3280
rect -3065 3250 -3055 3280
rect -3105 3240 -3055 3250
rect -3095 3075 -3055 3240
rect -3030 3230 -1835 3235
rect -3030 3195 -3020 3230
rect -1845 3195 -1835 3230
rect -3030 3175 -1835 3195
rect -3030 3140 -3020 3175
rect -1845 3140 -1835 3175
rect -3030 3120 -1835 3140
rect -3030 3085 -3020 3120
rect -1845 3085 -1835 3120
rect -3030 3080 -1835 3085
rect -3105 3065 -3055 3075
rect -3105 3035 -3095 3065
rect -3065 3035 -3055 3065
rect -3105 3025 -3055 3035
rect -3090 3020 -3055 3025
rect -3090 3015 -1835 3020
rect -3090 2985 -3020 3015
rect -1845 2985 -1835 3015
rect -3090 2980 -1835 2985
rect -2690 2915 -2650 2980
rect -3030 2905 -2980 2915
rect -3030 2875 -3020 2905
rect -2990 2875 -2980 2905
rect -3030 2865 -2980 2875
rect -2695 2905 -2645 2915
rect -2695 2875 -2685 2905
rect -2655 2875 -2645 2905
rect -2695 2865 -2645 2875
rect -1810 2905 -1760 2915
rect -1810 2875 -1800 2905
rect -1770 2875 -1760 2905
rect -1810 2865 -1760 2875
rect -3020 2845 -2990 2865
rect -1800 2845 -1770 2865
rect -3080 2835 -2985 2845
rect -3080 2830 -3020 2835
rect -3080 1665 -3070 2830
rect -3040 1665 -3020 2830
rect -3080 1660 -3020 1665
rect -2990 1660 -2985 2835
rect -3080 1645 -2985 1660
rect -2925 2835 -2875 2845
rect -2925 1660 -2920 2835
rect -2880 1660 -2875 2835
rect -2925 1615 -2875 1660
rect -2815 2835 -2775 2845
rect -2815 1660 -2810 2835
rect -2780 1660 -2775 2835
rect -2815 1650 -2775 1660
rect -2415 2835 -2375 2845
rect -2415 1660 -2410 2835
rect -2380 1660 -2375 2835
rect -3105 1570 -2875 1615
rect -3105 1535 -3070 1570
rect -2415 1535 -2375 1660
rect -2005 2835 -1965 2845
rect -2005 1660 -2000 2835
rect -1970 1660 -1965 2835
rect -2005 1650 -1965 1660
rect -1910 2835 -1860 2845
rect -1910 1660 -1900 2835
rect -1870 1660 -1860 2835
rect -1910 1615 -1860 1660
rect -1805 2835 -1710 2845
rect -1805 1660 -1800 2835
rect -1770 2830 -1710 2835
rect -1770 1665 -1750 2830
rect -1720 1665 -1710 2830
rect -1770 1660 -1710 1665
rect -1805 1645 -1710 1660
rect -1910 1570 -1675 1615
rect -1715 1535 -1675 1570
rect -3215 1525 -3165 1535
rect -3215 1495 -3205 1525
rect -3175 1495 -3165 1525
rect -3215 1485 -3165 1495
rect -3105 1525 -3015 1535
rect -3105 1495 -3055 1525
rect -3025 1495 -3015 1525
rect -3105 1485 -3015 1495
rect -2965 1525 -2915 1535
rect -2965 1495 -2955 1525
rect -2925 1520 -2915 1525
rect -2865 1525 -2815 1535
rect -2865 1520 -2855 1525
rect -2925 1495 -2855 1520
rect -2825 1520 -2815 1525
rect -2765 1525 -2715 1535
rect -2765 1520 -2755 1525
rect -2825 1495 -2755 1520
rect -2725 1520 -2715 1525
rect -2665 1525 -2615 1535
rect -2665 1520 -2655 1525
rect -2725 1495 -2655 1520
rect -2625 1520 -2615 1525
rect -2565 1525 -2215 1535
rect -2565 1520 -2555 1525
rect -2625 1495 -2555 1520
rect -2525 1500 -2455 1525
rect -2525 1495 -2515 1500
rect -2965 1485 -2515 1495
rect -2465 1495 -2455 1500
rect -2425 1500 -2355 1525
rect -2425 1495 -2415 1500
rect -2465 1485 -2415 1495
rect -2365 1495 -2355 1500
rect -2325 1500 -2255 1525
rect -2325 1495 -2315 1500
rect -2365 1485 -2315 1495
rect -2265 1495 -2255 1500
rect -2225 1520 -2215 1525
rect -2165 1525 -2115 1535
rect -2165 1520 -2155 1525
rect -2225 1495 -2155 1520
rect -2125 1520 -2115 1525
rect -2065 1525 -2015 1535
rect -2065 1520 -2055 1525
rect -2125 1495 -2055 1520
rect -2025 1520 -2015 1525
rect -1965 1525 -1915 1535
rect -1965 1520 -1955 1525
rect -2025 1495 -1955 1520
rect -1925 1520 -1915 1525
rect -1865 1525 -1815 1535
rect -1865 1520 -1855 1525
rect -1925 1495 -1855 1520
rect -1825 1495 -1815 1525
rect -2265 1485 -1815 1495
rect -1765 1525 -1675 1535
rect -1765 1495 -1755 1525
rect -1725 1495 -1675 1525
rect -1765 1485 -1675 1495
rect -1615 1525 -1565 1535
rect -1615 1495 -1605 1525
rect -1575 1495 -1565 1525
rect -1615 1485 -1565 1495
rect -3205 1465 -3175 1485
rect -3210 1455 -3170 1465
rect -3105 1460 -3070 1485
rect -3210 280 -3205 1455
rect -3175 280 -3170 1455
rect -3210 265 -3170 280
rect -3110 1455 -3070 1460
rect -3110 280 -3105 1455
rect -3075 280 -3070 1455
rect -3110 200 -3070 280
rect -3015 1455 -2965 1465
rect -3015 280 -3005 1455
rect -2975 280 -2965 1455
rect -3015 240 -2965 280
rect -2915 1455 -2865 1485
rect -2915 280 -2905 1455
rect -2875 280 -2865 1455
rect -2915 270 -2865 280
rect -2815 1455 -2765 1485
rect -2815 280 -2805 1455
rect -2775 280 -2765 1455
rect -2815 270 -2765 280
rect -2715 1455 -2665 1485
rect -2715 280 -2705 1455
rect -2675 280 -2665 1455
rect -2715 270 -2665 280
rect -2615 1455 -2565 1485
rect -2615 280 -2605 1455
rect -2575 280 -2565 1455
rect -2615 270 -2565 280
rect -2515 1455 -2465 1465
rect -2515 280 -2505 1455
rect -2475 280 -2465 1455
rect -2515 240 -2465 280
rect -2415 1455 -2365 1465
rect -2415 280 -2405 1455
rect -2375 280 -2365 1455
rect -2415 265 -2365 280
rect -2315 1455 -2265 1465
rect -2315 280 -2305 1455
rect -2275 280 -2265 1455
rect -2315 240 -2265 280
rect -2215 1455 -2165 1485
rect -2215 280 -2205 1455
rect -2175 280 -2165 1455
rect -2215 270 -2165 280
rect -2115 1455 -2065 1485
rect -2115 280 -2105 1455
rect -2075 280 -2065 1455
rect -2115 270 -2065 280
rect -2015 1455 -1965 1485
rect -2015 280 -2005 1455
rect -1975 280 -1965 1455
rect -2015 270 -1965 280
rect -1915 1455 -1865 1485
rect -1715 1470 -1675 1485
rect -1915 280 -1905 1455
rect -1875 280 -1865 1455
rect -1915 270 -1865 280
rect -1815 1455 -1765 1465
rect -1815 280 -1805 1455
rect -1775 280 -1765 1455
rect -1815 240 -1765 280
rect -1715 1455 -1665 1470
rect -1605 1465 -1575 1485
rect -1715 280 -1705 1455
rect -1675 280 -1665 1455
rect -1715 265 -1665 280
rect -1610 1455 -1570 1465
rect -1610 280 -1605 1455
rect -1575 280 -1570 1455
rect -1610 265 -1570 280
rect -3015 200 -1765 240
rect -1710 200 -1670 265
rect -3115 190 -3065 200
rect -3115 160 -3105 190
rect -3075 160 -3065 190
rect -1715 190 -1665 200
rect -1715 160 -1705 190
rect -1675 160 -1665 190
rect -3115 150 -1665 160
rect -3110 120 -1670 150
rect -2955 80 -1755 95
rect -2955 60 -2940 80
rect -1780 60 -1755 80
rect -2955 45 -1755 60
<< viali >>
rect -2980 7005 -1800 7035
rect -3205 5630 -3175 6805
rect -1605 5630 -1575 6805
rect -3010 4250 -2980 5425
rect -2810 4250 -2780 5425
rect -2000 4250 -1970 5425
rect -1800 4250 -1770 5425
rect -3020 3965 -1845 3995
rect -3020 3660 -1845 3690
rect -3020 3140 -1845 3175
rect -3020 1660 -2990 2835
rect -2810 1660 -2780 2835
rect -2000 1660 -1970 2835
rect -1800 1660 -1770 2835
rect -3205 280 -3175 1455
rect -2405 280 -2375 1455
rect -1605 280 -1575 1455
rect -2940 60 -1780 80
<< metal1 >>
rect -3215 7035 -1565 7040
rect -3215 7005 -2980 7035
rect -1800 7005 -1565 7035
rect -3215 6990 -1565 7005
rect -3215 6805 -3165 6990
rect -3215 5630 -3205 6805
rect -3175 5630 -3165 6805
rect -3215 2845 -3165 5630
rect -1615 6805 -1565 6990
rect -1615 5630 -1605 6805
rect -1575 5630 -1565 6805
rect -1615 5615 -1565 5630
rect -3020 5425 -2970 5440
rect -3020 4250 -3010 5425
rect -2980 4250 -2970 5425
rect -3020 4005 -2970 4250
rect -2820 5425 -2770 5440
rect -2820 4250 -2810 5425
rect -2780 4250 -2770 5425
rect -2820 4005 -2770 4250
rect -2010 5425 -1960 5445
rect -2010 4250 -2000 5425
rect -1970 4250 -1960 5425
rect -2010 4005 -1960 4250
rect -1810 5425 -1760 5440
rect -1810 4250 -1800 5425
rect -1770 4290 -1760 5425
rect -1770 4250 -1565 4290
rect -1810 4240 -1565 4250
rect -1615 4005 -1565 4240
rect -3030 3995 -1565 4005
rect -3030 3965 -3020 3995
rect -1845 3965 -1565 3995
rect -3030 3955 -1565 3965
rect -1615 3700 -1565 3955
rect -3030 3690 -1565 3700
rect -3030 3660 -3020 3690
rect -1845 3660 -1565 3690
rect -3030 3650 -1565 3660
rect -3030 3175 -1760 3185
rect -3030 3140 -3020 3175
rect -1845 3140 -1760 3175
rect -3030 3130 -1760 3140
rect -3215 2835 -2980 2845
rect -3215 2795 -3020 2835
rect -3030 1660 -3020 2795
rect -2990 1660 -2980 2835
rect -3030 1645 -2980 1660
rect -2820 2835 -2770 3130
rect -2820 1660 -2810 2835
rect -2780 1660 -2770 2835
rect -2820 1645 -2770 1660
rect -2010 2835 -1960 3130
rect -2010 1660 -2000 2835
rect -1970 1660 -1960 2835
rect -2010 1650 -1960 1660
rect -1810 2835 -1760 3130
rect -1810 1660 -1800 2835
rect -1770 1660 -1760 2835
rect -1810 1645 -1760 1660
rect -3215 1455 -3165 1470
rect -3215 280 -3205 1455
rect -3175 280 -3165 1455
rect -3215 105 -3165 280
rect -2415 1455 -2365 1470
rect -2415 280 -2405 1455
rect -2375 280 -2365 1455
rect -2415 105 -2365 280
rect -1615 1455 -1565 3650
rect -1615 280 -1605 1455
rect -1575 280 -1565 1455
rect -1615 105 -1565 280
rect -3215 80 -1565 105
rect -3215 60 -2940 80
rect -1780 60 -1565 80
rect -3215 55 -1565 60
<< end >>
