magic
tech sky130A
timestamp 1697752061
<< nwell >>
rect 1375 5485 3105 7030
<< poly >>
rect 1210 7370 1280 7400
rect 1250 7280 1280 7370
rect 1240 7270 1290 7280
rect 1240 7240 1250 7270
rect 1280 7240 1290 7270
rect 1240 7230 1290 7240
rect 1600 5455 1935 5475
rect 1600 4125 1650 5455
rect 1885 5415 1935 5455
rect 1480 4075 1650 4125
rect 1480 2905 1530 4075
rect 1320 2860 1530 2905
rect 1310 25 1360 35
rect 1310 -5 1320 25
rect 1350 -5 1360 25
rect 1310 -15 1360 -5
<< polycont >>
rect 1250 7240 1280 7270
rect 1320 -5 1350 25
<< locali >>
rect 1200 7300 1795 7330
rect 1240 7270 1290 7280
rect 1240 7240 1250 7270
rect 1280 7260 1290 7270
rect 1280 7240 1450 7260
rect 1240 7230 1450 7240
rect 1420 3805 1450 7230
rect 1765 6980 1795 7300
rect 1420 3775 1700 3805
rect 1660 3075 1695 3105
rect 1310 25 1360 35
rect 1310 -5 1320 25
rect 1350 10 1800 25
rect 1350 -5 1835 10
rect 1310 -15 1360 -5
use bias_generator  bias_generator_0
timestamp 1697739069
transform 1 0 4755 0 1 -45
box -3265 45 -1525 7075
use diffamp  diffamp_0
timestamp 1697750532
transform 1 0 750 0 1 6050
box -775 -6060 680 1350
<< labels >>
flabel space 1195 7365 1240 7395 0 FreeSans 168 0 0 0 Vbp
flabel locali 1210 7300 1255 7330 0 FreeSans 168 0 0 0 Vcp
flabel space 1305 2880 1350 2910 0 FreeSans 168 0 0 0 Vbn
flabel space 1260 5 1305 35 0 FreeSans 168 0 0 0 Vcn
flabel space 1325 4550 1375 4590 0 FreeSans 168 0 0 0 V1
flabel space 1390 3160 1440 3200 0 FreeSans 168 0 0 0 V2
<< end >>
