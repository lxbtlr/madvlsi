** LVS_BIASGEN flat netlist
*.OPIN VBP
*.OPIN VCN
*.OPIN VCP
*.OPIN VBN
*--------BEGIN_XM7->SKY130_FD_PR__PFET_01V8
XM7 VCP VDD VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM7->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM15->SKY130_FD_PR__PFET_01V8
XM15 VDD VDD NET2 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM15->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM16->SKY130_FD_PR__PFET_01V8
XM16 NET2 VDD NET1 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM16->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM17->SKY130_FD_PR__PFET_01V8
XM17 NET1 VDD VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM17->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM18->SKY130_FD_PR__PFET_01V8
XM18 VDD VDD NET5 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM18->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM19->SKY130_FD_PR__PFET_01V8
XM19 NET5 VDD VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM19->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM20->SKY130_FD_PR__PFET_01V8
XM20 VDD VDD NET3 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM20->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM21->SKY130_FD_PR__PFET_01V8
XM21 NET3 VDD NET4 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM21->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM22->SKY130_FD_PR__PFET_01V8
XM22 NET4 VDD VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM22->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM24->SKY130_FD_PR__PFET_01V8
XM24 VDD VDD VCP VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM24->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM25->SKY130_FD_PR__NFET_01V8
XM25 VCP VBN GND GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM25->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM14->SKY130_FD_PR__NFET_01V8
XM14 NET10 VBN GND GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM14->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM23->SKY130_FD_PR__NFET_01V8
XM23 NET11 VBN NET10 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM23->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM26->SKY130_FD_PR__NFET_01V8
XM26 NET12 VBN NET11 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM26->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM27->SKY130_FD_PR__NFET_01V8
XM27 NET13 VBN NET12 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM27->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM28->SKY130_FD_PR__NFET_01V8
XM28 VDD VBN NET13 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM28->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM29->SKY130_FD_PR__NFET_01V8
XM29 NET9 VBN VDD GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM29->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM30->SKY130_FD_PR__NFET_01V8
XM30 NET6 VBN NET9 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM30->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM31->SKY130_FD_PR__NFET_01V8
XM31 NET7 VBN NET6 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM31->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM32->SKY130_FD_PR__NFET_01V8
XM32 NET8 VBN NET7 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM32->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM33->SKY130_FD_PR__NFET_01V8
XM33 GND VBN NET8 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM33->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM34->SKY130_FD_PR__NFET_01V8
XM34 GND VBN VCP GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM34->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM35->SKY130_FD_PR__PFET_01V8
XM35 NET22 VBP VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM35->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM36->SKY130_FD_PR__PFET_01V8
XM36 VDD VBP NET16 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM36->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM37->SKY130_FD_PR__PFET_01V8
XM37 NET16 VBP NET14 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM37->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM38->SKY130_FD_PR__PFET_01V8
XM38 NET14 VBP NET15 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM38->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM39->SKY130_FD_PR__PFET_01V8
XM39 NET15 VBP NET20 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM39->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM40->SKY130_FD_PR__PFET_01V8
XM40 NET20 VBP NET17 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM40->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM41->SKY130_FD_PR__PFET_01V8
XM41 NET17 VBP NET18 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM41->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM42->SKY130_FD_PR__PFET_01V8
XM42 NET18 VBP NET19 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM42->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM43->SKY130_FD_PR__PFET_01V8
XM43 NET19 VBP VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM43->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM44->SKY130_FD_PR__PFET_01V8
XM44 VDD VBP NET21 VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM44->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM45->SKY130_FD_PR__NFET_01V8
XM45 VCN NET22 NET22 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM45->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM46->SKY130_FD_PR__NFET_01V8
XM46 NET20 NET20 NET23 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM46->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM47->SKY130_FD_PR__NFET_01V8
XM47 NET20 NET20 NET20 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM47->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM48->SKY130_FD_PR__NFET_01V8
XM48 NET20 NET20 NET20 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM48->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM49->SKY130_FD_PR__NFET_01V8
XM49 VCN NET20 NET20 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM49->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM50->SKY130_FD_PR__NFET_01V8
XM50 GND NET20 VCN GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM50->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM51->SKY130_FD_PR__NFET_01V8
XM51 VCN NET20 GND GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM51->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM52->SKY130_FD_PR__NFET_01V8
XM52 NET20 NET20 VCN GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM52->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM53->SKY130_FD_PR__NFET_01V8
XM53 NET20 NET20 NET20 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM53->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM54->SKY130_FD_PR__NFET_01V8
XM54 NET24 NET20 NET20 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM54->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM55->SKY130_FD_PR__NFET_01V8
XM55 NET20 NET20 NET24 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM55->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM56->SKY130_FD_PR__NFET_01V8
XM56 NET21 NET21 VCN GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM56->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM57->SKY130_FD_PR__NFET_01V8
XM57 GND VBN VBN GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM57->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM58->SKY130_FD_PR__NFET_01V8
XM58 VBP VBN GND GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM58->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM59->SKY130_FD_PR__PFET_01V8
XM59 VBP VBP VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM59->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM60->SKY130_FD_PR__NFET_01V8
XM60 GND VBN VBN GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM60->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM61->SKY130_FD_PR__NFET_01V8
XM61 VBP VBN GND GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM61->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM62->SKY130_FD_PR__PFET_01V8
XM62 VBP VBP VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM62->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM1->SKY130_FD_PR__PFET_01V8
XM1 NET21 VDD VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM1->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM2->SKY130_FD_PR__NFET_01V8
XM2 GND GND NET21 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM2->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM3->SKY130_FD_PR__PFET_01V8
XM3 NET22 VDD VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM3->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM4->SKY130_FD_PR__NFET_01V8
XM4 GND GND NET22 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM4->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM5->SKY130_FD_PR__PFET_01V8
XM5 VCP VDD VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM5->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM6->SKY130_FD_PR__NFET_01V8
XM6 GND GND VCP GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM6->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM8->SKY130_FD_PR__PFET_01V8
XM8 VCP VDD VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM8->SKY130_FD_PR__PFET_01V8
*--------BEGIN_XM9->SKY130_FD_PR__NFET_01V8
XM9 GND GND VCP GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM9->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM10->SKY130_FD_PR__NFET_01V8
XM10 VCN NET20 NET20 GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM10->SKY130_FD_PR__NFET_01V8
*--------BEGIN_XM11->SKY130_FD_PR__NFET_01V8
XM11 NET23 NET20 VCN GND  SKY130_FD_PR__NFET_01V8 L=0.5 W=12 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29'
+ PD='2*INT((NF+1)/2)*(W/NF+0.29)' PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0
+ SD=0 MULT=1 M=1
*--------END___XM11->SKY130_FD_PR__NFET_01V8
.end
