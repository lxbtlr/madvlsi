magic
tech sky130A
timestamp 1695856067
<< nwell >>
rect -115 620 345 1165
<< nmos >>
rect -65 445 -50 545
rect 0 445 15 545
rect -10 245 5 345
rect 210 345 225 545
rect 250 345 265 545
rect -10 95 5 195
rect 180 95 195 195
rect 245 95 260 195
<< pmos >>
rect 5 1005 20 1105
rect 70 1005 85 1105
rect 220 945 235 1145
rect 260 945 275 1145
rect -25 830 -10 930
rect -25 670 -10 770
rect 185 645 200 745
rect 250 645 265 745
<< ndiff >>
rect -115 530 -65 545
rect -115 460 -100 530
rect -80 460 -65 530
rect -115 445 -65 460
rect -50 530 0 545
rect -50 460 -35 530
rect -15 460 0 530
rect -50 445 0 460
rect 15 530 65 545
rect 15 460 30 530
rect 50 460 65 530
rect 15 445 65 460
rect 160 530 210 545
rect -60 330 -10 345
rect -60 260 -45 330
rect -25 260 -10 330
rect -60 245 -10 260
rect 5 330 55 345
rect 5 260 20 330
rect 40 260 55 330
rect 5 245 55 260
rect 160 360 175 530
rect 195 360 210 530
rect 160 345 210 360
rect 225 345 250 545
rect 265 530 315 545
rect 265 360 280 530
rect 300 360 315 530
rect 265 345 315 360
rect -60 180 -10 195
rect -60 110 -45 180
rect -25 110 -10 180
rect -60 95 -10 110
rect 5 180 55 195
rect 5 110 20 180
rect 40 110 55 180
rect 5 95 55 110
rect 135 180 180 195
rect 135 110 145 180
rect 165 110 180 180
rect 135 95 180 110
rect 195 180 245 195
rect 195 110 210 180
rect 230 110 245 180
rect 195 95 245 110
rect 260 180 310 195
rect 260 110 275 180
rect 295 110 310 180
rect 260 95 310 110
<< pdiff >>
rect 170 1130 220 1145
rect -44 1090 5 1105
rect -44 1020 -30 1090
rect -10 1020 5 1090
rect -44 1005 5 1020
rect 20 1090 70 1105
rect 20 1020 35 1090
rect 55 1020 70 1090
rect 20 1005 70 1020
rect 85 1090 135 1105
rect 85 1020 100 1090
rect 120 1020 135 1090
rect 85 1005 135 1020
rect 170 960 185 1130
rect 205 960 220 1130
rect 170 945 220 960
rect 235 945 260 1145
rect 275 1130 325 1145
rect 275 960 290 1130
rect 310 960 325 1130
rect 275 945 325 960
rect -75 915 -25 930
rect -75 845 -60 915
rect -40 845 -25 915
rect -75 830 -25 845
rect -10 915 40 930
rect -10 845 5 915
rect 25 845 40 915
rect -10 830 40 845
rect -75 755 -25 770
rect -75 685 -60 755
rect -40 685 -25 755
rect -75 670 -25 685
rect -10 755 40 770
rect -10 685 5 755
rect 25 685 40 755
rect -10 670 40 685
rect 140 730 185 745
rect 140 660 150 730
rect 170 660 185 730
rect 140 645 185 660
rect 200 730 250 745
rect 200 660 215 730
rect 235 660 250 730
rect 200 645 250 660
rect 265 730 315 745
rect 265 660 280 730
rect 300 660 315 730
rect 265 645 315 660
<< ndiffc >>
rect -100 460 -80 530
rect -35 460 -15 530
rect 30 460 50 530
rect -45 260 -25 330
rect 20 260 40 330
rect 175 360 195 530
rect 280 360 300 530
rect -45 110 -25 180
rect 20 110 40 180
rect 145 110 165 180
rect 210 110 230 180
rect 275 110 295 180
<< pdiffc >>
rect -30 1020 -10 1090
rect 35 1020 55 1090
rect 100 1020 120 1090
rect 185 960 205 1130
rect 290 960 310 1130
rect -60 845 -40 915
rect 5 845 25 915
rect -60 685 -40 755
rect 5 685 25 755
rect 150 660 170 730
rect 215 660 235 730
rect 280 660 300 730
<< psubdiff >>
rect -110 180 -60 195
rect -110 110 -95 180
rect -75 110 -60 180
rect -110 95 -60 110
<< psubdiffcont >>
rect -95 110 -75 180
<< poly >>
rect -85 1160 -40 1165
rect -85 1155 85 1160
rect -85 1130 -75 1155
rect -50 1145 85 1155
rect 220 1145 235 1160
rect 260 1145 275 1160
rect -50 1130 -40 1145
rect -85 1120 -40 1130
rect 5 1105 20 1120
rect 70 1105 85 1145
rect 5 990 20 1005
rect 70 990 85 1005
rect -100 980 -55 990
rect -100 955 -90 980
rect -65 955 -55 980
rect 5 975 40 990
rect -100 945 -55 955
rect 25 965 40 975
rect 25 955 135 965
rect 25 950 100 955
rect -100 630 -85 945
rect -25 930 -10 945
rect 90 930 100 950
rect 125 930 135 955
rect 90 920 135 930
rect 220 925 235 945
rect 260 925 275 945
rect 160 910 275 925
rect 160 895 175 910
rect 75 880 175 895
rect -25 815 -10 830
rect 75 815 90 880
rect -25 800 90 815
rect 155 835 200 845
rect 155 810 165 835
rect 190 810 200 835
rect 155 800 200 810
rect 285 840 330 850
rect 285 815 295 840
rect 320 815 330 840
rect 285 805 330 815
rect -25 770 -10 800
rect 185 745 200 800
rect 300 775 315 805
rect 250 760 315 775
rect 250 745 265 760
rect -25 655 -10 670
rect -25 640 65 655
rect -100 620 -55 630
rect -100 595 -90 620
rect -65 600 -55 620
rect -65 595 15 600
rect -100 585 15 595
rect -65 545 -50 560
rect 0 545 15 585
rect 50 570 65 640
rect 185 630 200 645
rect 120 610 165 620
rect 120 585 130 610
rect 155 605 165 610
rect 250 605 265 645
rect 155 590 265 605
rect 155 585 165 590
rect 120 575 165 585
rect 50 555 95 570
rect 80 455 95 555
rect 210 545 225 560
rect 250 545 265 560
rect -65 405 -50 445
rect 0 430 15 445
rect 80 440 115 455
rect 30 405 75 410
rect -65 400 75 405
rect -65 390 40 400
rect 30 375 40 390
rect 65 375 75 400
rect 30 365 75 375
rect -10 345 5 360
rect 100 335 115 440
rect 210 335 225 345
rect 250 335 265 345
rect 100 320 265 335
rect -10 225 5 245
rect 100 225 115 320
rect 165 285 210 295
rect 165 260 175 285
rect 200 260 210 285
rect 165 250 210 260
rect -10 210 115 225
rect -10 195 5 210
rect 180 195 195 250
rect 235 245 280 255
rect 235 220 245 245
rect 270 220 280 245
rect 235 210 280 220
rect 245 195 260 210
rect -10 80 5 95
rect 180 80 195 95
rect 245 80 260 95
<< polycont >>
rect -75 1130 -50 1155
rect -90 955 -65 980
rect 100 930 125 955
rect 165 810 190 835
rect 295 815 320 840
rect -90 595 -65 620
rect 130 585 155 610
rect 40 375 65 400
rect 175 260 200 285
rect 245 220 270 245
<< locali >>
rect -85 1155 -40 1165
rect -85 1130 -75 1155
rect -50 1130 -40 1155
rect -85 1120 -40 1130
rect -60 1100 -40 1120
rect 175 1130 215 1140
rect -60 1090 0 1100
rect -60 1020 -30 1090
rect -10 1020 0 1090
rect -60 1010 0 1020
rect 25 1090 65 1100
rect 25 1020 35 1090
rect 55 1020 65 1090
rect 25 1010 65 1020
rect 90 1090 130 1100
rect 90 1020 100 1090
rect 120 1020 130 1090
rect 90 1010 130 1020
rect -60 1002 -40 1010
rect -77 990 -40 1002
rect -100 980 -40 990
rect -100 955 -90 980
rect -65 955 -55 980
rect 105 965 125 1010
rect -100 945 -55 955
rect 90 955 135 965
rect 90 945 100 955
rect 15 930 100 945
rect 125 930 135 955
rect 15 925 135 930
rect -70 915 -30 925
rect -70 890 -60 915
rect -115 870 -60 890
rect -70 845 -60 870
rect -40 845 -30 915
rect -70 835 -30 845
rect -5 915 35 925
rect 90 920 135 925
rect 175 960 185 1130
rect 205 960 215 1130
rect 175 955 215 960
rect 280 1130 320 1140
rect 280 960 290 1130
rect 310 960 320 1130
rect -5 845 5 915
rect 25 855 35 915
rect 175 900 195 955
rect 280 950 320 960
rect 115 880 195 900
rect 25 845 75 855
rect -5 835 75 845
rect -115 765 -45 780
rect -115 760 -30 765
rect -70 755 -30 760
rect -70 685 -60 755
rect -40 685 -30 755
rect -70 675 -30 685
rect -5 755 35 765
rect -5 685 5 755
rect 25 685 35 755
rect -5 675 35 685
rect -5 655 15 675
rect -25 635 15 655
rect -100 620 -55 630
rect -25 620 -5 635
rect 55 620 75 835
rect 115 780 135 880
rect 245 870 340 890
rect 155 835 200 845
rect 155 810 165 835
rect 190 825 200 835
rect 245 825 265 870
rect 190 810 265 825
rect 155 805 265 810
rect 285 840 330 850
rect 285 815 295 840
rect 320 815 330 840
rect 285 805 330 815
rect 155 800 200 805
rect 245 785 265 805
rect 115 760 225 780
rect 245 765 290 785
rect 205 740 225 760
rect 270 740 290 765
rect 310 780 330 805
rect 310 760 340 780
rect 140 730 180 740
rect 140 660 150 730
rect 170 660 180 730
rect 140 650 180 660
rect 205 730 245 740
rect 205 660 215 730
rect 235 660 245 730
rect 205 650 245 660
rect 270 730 310 740
rect 270 660 280 730
rect 300 660 310 730
rect 270 650 310 660
rect 140 620 160 650
rect -100 595 -90 620
rect -65 600 -5 620
rect 25 600 75 620
rect 120 610 165 620
rect -65 595 -55 600
rect -100 585 -55 595
rect -100 540 -80 585
rect 25 540 45 600
rect 120 585 130 610
rect 155 585 165 610
rect 120 575 165 585
rect -110 530 -70 540
rect -110 460 -100 530
rect -80 460 -70 530
rect -110 450 -70 460
rect -45 530 -5 540
rect -45 460 -35 530
rect -15 460 -5 530
rect -45 450 -5 460
rect 20 530 60 540
rect 20 460 30 530
rect 50 460 60 530
rect 20 450 60 460
rect -45 430 -25 450
rect -95 410 -25 430
rect 30 410 50 450
rect -95 190 -75 410
rect 30 400 75 410
rect 30 385 40 400
rect -35 375 40 385
rect 65 375 75 400
rect -35 365 75 375
rect -35 340 -15 365
rect -55 330 -15 340
rect -55 260 -45 330
rect -25 260 -15 330
rect -55 250 -15 260
rect 10 330 50 340
rect 10 260 20 330
rect 40 270 50 330
rect 125 270 145 575
rect 275 540 295 650
rect 165 530 205 540
rect 165 360 175 530
rect 195 360 205 530
rect 165 350 205 360
rect 270 530 310 540
rect 270 360 280 530
rect 300 360 310 530
rect 270 350 310 360
rect 290 295 310 350
rect 40 260 145 270
rect 10 250 145 260
rect 165 285 320 295
rect 165 260 175 285
rect 200 275 320 285
rect 200 260 210 275
rect 165 250 210 260
rect 125 230 145 250
rect 235 245 280 255
rect 235 230 245 245
rect 125 220 245 230
rect 270 220 280 245
rect 125 210 280 220
rect 135 190 152 210
rect 300 190 320 275
rect -105 180 -15 190
rect -105 110 -95 180
rect -75 110 -45 180
rect -25 110 -15 180
rect -105 100 -15 110
rect 10 180 55 190
rect 10 110 20 180
rect 40 110 55 180
rect 10 100 55 110
rect 135 180 175 190
rect 135 110 145 180
rect 165 110 175 180
rect 135 100 175 110
rect 200 180 240 190
rect 200 110 210 180
rect 230 110 240 180
rect 200 100 240 110
rect 265 180 320 190
rect 265 110 275 180
rect 295 165 320 180
rect 295 110 305 165
rect 265 100 305 110
<< viali >>
rect 35 1020 55 1090
rect 290 960 310 1130
rect -100 460 -80 530
rect 175 360 195 530
rect 20 110 40 180
rect 210 110 230 180
<< metal1 >>
rect -115 1130 340 1155
rect -115 1090 290 1130
rect -115 1020 35 1090
rect 55 1020 290 1090
rect -115 960 290 1020
rect 310 960 340 1130
rect -115 950 340 960
rect -115 530 340 545
rect -115 460 -100 530
rect -80 460 175 530
rect -115 360 175 460
rect 195 360 340 530
rect -115 345 340 360
rect -115 180 340 195
rect -115 110 20 180
rect 40 110 210 180
rect 230 110 340 180
rect -115 95 340 110
<< labels >>
rlabel metal1 -115 400 -115 400 7 CLK
port 5 w
rlabel metal1 -115 140 -115 140 7 VN
port 6 w
rlabel metal1 -115 1040 -115 1040 7 VP
port 7 w
rlabel locali -115 770 -115 770 7 D
port 2 w
rlabel locali -115 880 -115 880 7 D_NOT
port 1 w
rlabel locali 340 770 340 770 7 Q_NOT
port 3 w
rlabel locali 340 880 340 880 7 Q
port 4 w
<< end >>
